
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_windowed_RF is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_windowed_RF;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_RF.all;

entity register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_4 is

   port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (4 downto 0);  CO : out std_logic);

end register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_4;

architecture SYN_rpl of register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, carry_2_port, carry_1_port, n1 : 
      std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => n1, S
                           => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => carry_1_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_RF.all;

entity register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_3 is

   port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (4 downto 0);  CO : out std_logic);

end register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_3;

architecture SYN_rpl of register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, carry_2_port, carry_1_port, n1 : 
      std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => n1, S
                           => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => carry_1_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_RF.all;

entity register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_2 is

   port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (4 downto 0);  CO : out std_logic);

end register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_2;

architecture SYN_rpl of register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, carry_2_port, carry_1_port, n1 : 
      std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => n1, S
                           => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => carry_1_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_RF.all;

entity register_CU_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_incdec_0 is

   port( A : in std_logic_vector (4 downto 0);  INC_DEC : in std_logic;  SUM : 
         out std_logic_vector (4 downto 0));

end register_CU_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_incdec_0;

architecture SYN_rpl of register_CU_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_incdec_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, carry_2_port, carry_1_port, carry_0_port,
      n1 : std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => INC_DEC, CI => carry_4_port, CO => n1
                           , S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => INC_DEC, CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => INC_DEC, CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => INC_DEC, CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => INC_DEC, CI => carry_0_port, CO => 
                           carry_1_port, S => SUM(0));
   U1 : INV_X1 port map( A => INC_DEC, ZN => carry_0_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_RF.all;

entity register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3 is

   port( clk, reset, enable, call, ret : in std_logic;  datain : in 
         std_logic_vector (63 downto 0);  rd1, rd2, wr : in std_logic;  add_wr,
         add_rd1, add_rd2 : in std_logic_vector (4 downto 0);  in_from_mem : in
         std_logic_vector (63 downto 0);  cwp : in std_logic_vector (1 downto 
         0);  count3 : in std_logic_vector (3 downto 0);  spill, fill : in 
         std_logic;  out_to_mem, out1, out2 : out std_logic_vector (63 downto 
         0));

end register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3;

architecture SYN_bhv of register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_4
      port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (4 downto 0);  CO : out std_logic);
   end component;
   
   component register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_3
      port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (4 downto 0);  CO : out std_logic);
   end component;
   
   component register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_2
      port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (4 downto 0);  CO : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal out_to_mem_63_port, out_to_mem_62_port, out_to_mem_61_port, 
      out_to_mem_60_port, out_to_mem_59_port, out_to_mem_58_port, 
      out_to_mem_57_port, out_to_mem_56_port, out_to_mem_55_port, 
      out_to_mem_54_port, out_to_mem_53_port, out_to_mem_52_port, 
      out_to_mem_51_port, out_to_mem_50_port, out_to_mem_49_port, 
      out_to_mem_48_port, out_to_mem_47_port, out_to_mem_46_port, 
      out_to_mem_45_port, out_to_mem_44_port, out_to_mem_43_port, 
      out_to_mem_42_port, out_to_mem_41_port, out_to_mem_40_port, 
      out_to_mem_39_port, out_to_mem_38_port, out_to_mem_37_port, 
      out_to_mem_36_port, out_to_mem_35_port, out_to_mem_34_port, 
      out_to_mem_33_port, out_to_mem_32_port, out_to_mem_31_port, 
      out_to_mem_30_port, out_to_mem_29_port, out_to_mem_28_port, 
      out_to_mem_27_port, out_to_mem_26_port, out_to_mem_25_port, 
      out_to_mem_24_port, out_to_mem_23_port, out_to_mem_22_port, 
      out_to_mem_21_port, out_to_mem_20_port, out_to_mem_19_port, 
      out_to_mem_18_port, out_to_mem_17_port, out_to_mem_16_port, 
      out_to_mem_15_port, out_to_mem_14_port, out_to_mem_13_port, 
      out_to_mem_12_port, out_to_mem_11_port, out_to_mem_10_port, 
      out_to_mem_9_port, out_to_mem_8_port, out_to_mem_7_port, 
      out_to_mem_6_port, out_to_mem_5_port, out_to_mem_4_port, 
      out_to_mem_3_port, out_to_mem_2_port, out_to_mem_1_port, 
      out_to_mem_0_port, N78, N79, N80, N92, N113, N114, N115, N127, N148, N149
      , N150, N162, registers_15_63_port, registers_15_62_port, 
      registers_15_61_port, registers_15_60_port, registers_15_59_port, 
      registers_15_58_port, registers_15_57_port, registers_15_56_port, 
      registers_15_55_port, registers_15_54_port, registers_15_53_port, 
      registers_15_52_port, registers_15_51_port, registers_15_50_port, 
      registers_15_49_port, registers_15_48_port, registers_15_47_port, 
      registers_15_46_port, registers_15_45_port, registers_15_44_port, 
      registers_15_43_port, registers_15_42_port, registers_15_41_port, 
      registers_15_40_port, registers_15_39_port, registers_15_38_port, 
      registers_15_37_port, registers_15_36_port, registers_15_35_port, 
      registers_15_34_port, registers_15_33_port, registers_15_32_port, 
      registers_15_31_port, registers_15_30_port, registers_15_29_port, 
      registers_15_28_port, registers_15_27_port, registers_15_26_port, 
      registers_15_25_port, registers_15_24_port, registers_15_23_port, 
      registers_15_22_port, registers_15_21_port, registers_15_20_port, 
      registers_15_19_port, registers_15_18_port, registers_15_17_port, 
      registers_15_16_port, registers_15_15_port, registers_15_14_port, 
      registers_15_13_port, registers_15_12_port, registers_15_11_port, 
      registers_15_10_port, registers_15_9_port, registers_15_8_port, 
      registers_15_7_port, registers_15_6_port, registers_15_5_port, 
      registers_15_4_port, registers_15_3_port, registers_15_2_port, 
      registers_15_1_port, registers_15_0_port, registers_14_63_port, 
      registers_14_62_port, registers_14_61_port, registers_14_60_port, 
      registers_14_59_port, registers_14_58_port, registers_14_57_port, 
      registers_14_56_port, registers_14_55_port, registers_14_54_port, 
      registers_14_53_port, registers_14_52_port, registers_14_51_port, 
      registers_14_50_port, registers_14_49_port, registers_14_48_port, 
      registers_14_47_port, registers_14_46_port, registers_14_45_port, 
      registers_14_44_port, registers_14_43_port, registers_14_42_port, 
      registers_14_41_port, registers_14_40_port, registers_14_39_port, 
      registers_14_38_port, registers_14_37_port, registers_14_36_port, 
      registers_14_35_port, registers_14_34_port, registers_14_33_port, 
      registers_14_32_port, registers_14_31_port, registers_14_30_port, 
      registers_14_29_port, registers_14_28_port, registers_14_27_port, 
      registers_14_26_port, registers_14_25_port, registers_14_24_port, 
      registers_14_23_port, registers_14_22_port, registers_14_21_port, 
      registers_14_20_port, registers_14_19_port, registers_14_18_port, 
      registers_14_17_port, registers_14_16_port, registers_14_15_port, 
      registers_14_14_port, registers_14_13_port, registers_14_12_port, 
      registers_14_11_port, registers_14_10_port, registers_14_9_port, 
      registers_14_8_port, registers_14_7_port, registers_14_6_port, 
      registers_14_5_port, registers_14_4_port, registers_14_3_port, 
      registers_14_2_port, registers_14_1_port, registers_14_0_port, 
      registers_4_63_port, registers_4_62_port, registers_4_61_port, 
      registers_4_60_port, registers_4_59_port, registers_4_58_port, 
      registers_4_57_port, registers_4_56_port, registers_4_55_port, 
      registers_4_54_port, registers_4_53_port, registers_4_52_port, 
      registers_4_51_port, registers_4_50_port, registers_4_49_port, 
      registers_4_48_port, registers_4_47_port, registers_4_46_port, 
      registers_4_45_port, registers_4_44_port, registers_4_43_port, 
      registers_4_42_port, registers_4_41_port, registers_4_40_port, 
      registers_4_39_port, registers_4_38_port, registers_4_37_port, 
      registers_4_36_port, registers_4_35_port, registers_4_34_port, 
      registers_4_33_port, registers_4_32_port, registers_4_31_port, 
      registers_4_30_port, registers_4_29_port, registers_4_28_port, 
      registers_4_27_port, registers_4_26_port, registers_4_25_port, 
      registers_4_24_port, registers_4_23_port, registers_4_22_port, 
      registers_4_21_port, registers_4_20_port, registers_4_19_port, 
      registers_4_18_port, registers_4_17_port, registers_4_16_port, 
      registers_4_15_port, registers_4_14_port, registers_4_13_port, 
      registers_4_12_port, registers_4_11_port, registers_4_10_port, 
      registers_4_9_port, registers_4_8_port, registers_4_7_port, 
      registers_4_6_port, registers_4_5_port, registers_4_4_port, 
      registers_4_3_port, registers_4_2_port, registers_4_1_port, 
      registers_4_0_port, registers_3_63_port, registers_3_62_port, 
      registers_3_61_port, registers_3_60_port, registers_3_59_port, 
      registers_3_58_port, registers_3_57_port, registers_3_56_port, 
      registers_3_55_port, registers_3_54_port, registers_3_53_port, 
      registers_3_52_port, registers_3_51_port, registers_3_50_port, 
      registers_3_49_port, registers_3_48_port, registers_3_47_port, 
      registers_3_46_port, registers_3_45_port, registers_3_44_port, 
      registers_3_43_port, registers_3_42_port, registers_3_41_port, 
      registers_3_40_port, registers_3_39_port, registers_3_38_port, 
      registers_3_37_port, registers_3_36_port, registers_3_35_port, 
      registers_3_34_port, registers_3_33_port, registers_3_32_port, 
      registers_3_31_port, registers_3_30_port, registers_3_29_port, 
      registers_3_28_port, registers_3_27_port, registers_3_26_port, 
      registers_3_25_port, registers_3_24_port, registers_3_23_port, 
      registers_3_22_port, registers_3_21_port, registers_3_20_port, 
      registers_3_19_port, registers_3_18_port, registers_3_17_port, 
      registers_3_16_port, registers_3_15_port, registers_3_14_port, 
      registers_3_13_port, registers_3_12_port, registers_3_11_port, 
      registers_3_10_port, registers_3_9_port, registers_3_8_port, 
      registers_3_7_port, registers_3_6_port, registers_3_5_port, 
      registers_3_4_port, registers_3_3_port, registers_3_2_port, 
      registers_3_1_port, registers_3_0_port, U3_U2_Z_0, U3_U2_Z_1, U3_U2_Z_2, 
      U3_U2_Z_3, U3_U2_Z_4, U3_U4_Z_0, U3_U4_Z_1, U3_U4_Z_2, U3_U4_Z_3, 
      U3_U4_Z_4, U3_U6_Z_0, U3_U6_Z_1, U3_U6_Z_2, U3_U6_Z_3, U3_U6_Z_4, n7023, 
      n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, 
      n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, 
      n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, 
      n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, 
      n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, 
      n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, 
      n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, 
      n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, 
      n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, 
      n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, 
      n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, 
      n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, 
      n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, 
      n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, 
      n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, 
      n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, 
      n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, 
      n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, 
      n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, 
      n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, 
      n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, 
      n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, 
      n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, 
      n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, 
      n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, 
      n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, 
      n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, 
      n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, 
      n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, 
      n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, 
      n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, 
      n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, 
      n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, 
      n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, 
      n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, 
      n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, 
      n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, 
      n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, 
      n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, 
      n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, 
      n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, 
      n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, 
      n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, 
      n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, 
      n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, 
      n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, 
      n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, 
      n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, 
      n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, 
      n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, 
      n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, 
      n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, 
      n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, 
      n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, 
      n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, 
      n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, 
      n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, 
      n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, 
      n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, 
      n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, 
      n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, 
      n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, 
      n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, 
      n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, 
      n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, 
      n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, 
      n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, 
      n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, 
      n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, 
      n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, 
      n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, 
      n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, 
      n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, 
      n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, 
      n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, 
      n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, 
      n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, 
      n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, 
      n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, 
      n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, 
      n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, 
      n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, 
      n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, 
      n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, 
      n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, 
      n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, 
      n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, 
      n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, 
      n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, 
      n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, 
      n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, 
      n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, 
      n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, 
      n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, 
      n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, 
      n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, 
      n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, 
      n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, 
      n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, 
      n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, 
      n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, 
      n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, 
      n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, 
      n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, 
      n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, 
      n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, 
      n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, 
      n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, 
      n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, 
      n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, 
      n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, 
      n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, 
      n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, 
      n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, 
      n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, 
      n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, 
      n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, 
      n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, 
      n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, 
      n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, 
      n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, 
      n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, 
      n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, 
      n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, 
      n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, 
      n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, 
      n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, 
      n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, 
      n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, 
      n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, 
      n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, 
      n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, 
      n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, 
      n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, 
      n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, 
      n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, 
      n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, 
      n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, 
      n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, 
      n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, 
      n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, 
      n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, 
      n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, 
      n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, 
      n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, 
      n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, 
      n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, 
      n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, 
      n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, 
      n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, 
      n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, 
      n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, 
      n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, 
      n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, 
      n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, 
      n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, 
      n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, 
      n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, 
      n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, 
      n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, 
      n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, 
      n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, 
      n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, 
      n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, 
      n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, 
      n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, 
      n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, 
      n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, 
      n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, 
      n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, 
      n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, 
      n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, 
      n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, 
      n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, 
      n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, 
      n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, 
      n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, 
      n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, 
      n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, 
      n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, 
      n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, 
      n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, 
      n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, 
      n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, 
      n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, 
      n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, 
      n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, 
      n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, 
      n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, 
      n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, 
      n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, 
      n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, 
      n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, 
      n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, 
      n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, 
      n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, 
      n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, 
      n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, 
      n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, 
      n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, 
      n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, 
      n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, 
      n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, 
      n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, 
      n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, 
      n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, 
      n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, 
      n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, 
      n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, 
      n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, 
      n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, 
      n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, 
      n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, 
      n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, 
      n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, 
      n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, 
      n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, 
      n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, 
      n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, 
      n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, 
      n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, 
      n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, 
      n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, 
      n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, 
      sub_105_carry_4_port, sub_86_carry_4_port, sub_123_carry_4_port, n2145, 
      n2146, n2148, n2149, n2151, n2152, n2154, n2155, n2157, n2158, n2160, 
      n2161, n2163, n2164, n2166, n2167, n2169, n2170, n2172, n2173, n2175, 
      n2176, n2178, n2179, n2181, n2182, n2184, n2185, n2187, n2188, n2190, 
      n2191, n2193, n2194, n2196, n2197, n2199, n2200, n2202, n2203, n2205, 
      n2206, n2208, n2209, n2211, n2212, n2214, n2215, n2217, n2218, n2220, 
      n2221, n2223, n2224, n2226, n2227, n2229, n2230, n2232, n2233, n2235, 
      n2236, n2238, n2239, n2241, n2242, n2244, n2245, n2247, n2248, n2250, 
      n2251, n2253, n2254, n2256, n2257, n2259, n2260, n2262, n2263, n2265, 
      n2266, n2268, n2269, n2271, n2272, n2274, n2275, n2277, n2278, n2280, 
      n2281, n2283, n2284, n2286, n2287, n2289, n2290, n2292, n2293, n2295, 
      n2296, n2298, n2299, n2301, n2302, n2304, n2305, n2307, n2308, n2310, 
      n2311, n2313, n2314, n2316, n2317, n2319, n2320, n2322, n2323, n2325, 
      n2326, n2328, n2329, n2331, n2332, n2334, n2335, n3169, n3171, n3173, 
      n3175, n3177, n3179, n3181, n3183, n3185, n3187, n3189, n3191, n3193, 
      n3195, n3197, n3199, n3201, n3203, n3205, n3207, n3209, n3211, n3213, 
      n3215, n3217, n3219, n3221, n3223, n3225, n3227, n3229, n3231, n3233, 
      n3235, n3237, n3239, n3241, n3243, n3245, n3247, n3249, n3251, n3253, 
      n3255, n3257, n3259, n3261, n3263, n3265, n3267, n3269, n3271, n3273, 
      n3275, n3277, n3279, n3281, n3283, n3285, n3287, n3289, n3291, n3293, 
      n3295, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, 
      n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, 
      n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, 
      n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, 
      n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, 
      n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, 
      n3362, n3363, n3364, n3365, n3366, n3371, n3372, n3373, n3374, n3375, 
      n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, 
      n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, 
      n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, 
      n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, 
      n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, 
      n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3439, 
      n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, 
      n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, 
      n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, 
      n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, 
      n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, 
      n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, 
      n3500, n3501, n3502, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
      n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, 
      n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, 
      n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, 
      n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, 
      n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, 
      n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3574, n3575, n3576, 
      n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, 
      n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, 
      n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, 
      n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, 
      n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, 
      n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, 
      n3637, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, 
      n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, 
      n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, 
      n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, 
      n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, 
      n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, 
      n3700, n3701, n3702, n3703, n3704, n3707, n3708, n3709, n3710, n3711, 
      n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, 
      n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, 
      n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, 
      n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, 
      n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, 
      n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3773, 
      n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, 
      n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, 
      n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, 
      n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, 
      n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, 
      n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, 
      n3834, n3835, n3836, n3974, n3975, n3976, n3977, n3978, n3979, n3980, 
      n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, 
      n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, 
      n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, 
      n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, 
      n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, 
      n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4040, n4041, n4042, 
      n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, 
      n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, 
      n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, 
      n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, 
      n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, 
      n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, 
      n4103, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, 
      n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, 
      n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, 
      n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, 
      n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, 
      n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, 
      n4238, n4239, n4240, n4241, n4242, n4246, n4247, n4248, n4249, n4250, 
      n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, 
      n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, 
      n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, 
      n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, 
      n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, 
      n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4448, 
      n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, 
      n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, 
      n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, 
      n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, 
      n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, 
      n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, 
      n4509, n4510, n4511, n4517, n4518, n4519, n4520, n4521, n4522, n4523, 
      n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, 
      n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, 
      n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, 
      n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, 
      n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, 
      n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4654, n4655, n4656, 
      n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, 
      n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, 
      n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, 
      n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, 
      n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, 
      n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, 
      n4717, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, 
      n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, 
      n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, 
      n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, 
      n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, 
      n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, 
      n4779, n4780, n4781, n4782, n4783, n4787, n4788, n4789, n4790, n4791, 
      n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, 
      n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, 
      n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, 
      n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, 
      n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, 
      n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4858, 
      n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, 
      n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, 
      n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, 
      n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, 
      n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, 
      n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, 
      n4919, n4920, n4921, n4924, n4925, n4926, n4927, n4928, n4929, n4930, 
      n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, 
      n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, 
      n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, 
      n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, 
      n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, 
      n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4990, n4991, n4992, 
      n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, 
      n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, 
      n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, 
      n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, 
      n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, 
      n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, 
      n5053, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, 
      n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, 
      n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, 
      n5286, n5287, n5288, n5289, n5290, n5291, n5355, n5356, n5357, n5359, 
      n5424, n5426, n5491, n5492, n5494, n5559, n5560, n5562, n5627, n5629, 
      n5694, n5695, n5696, n5698, n5763, n5764, n5765, n5766, n5767, n5769, 
      n5835, n5901, n5966, n5968, n6033, n15077, n15078, n15079, n15297, n15298
      , n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
      n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, 
      n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, 
      n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, 
      n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, 
      n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, 
      n15353, n15354, n15355, n15356, n15417, n15418, n15419, n15420, n15421, 
      n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, 
      n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, 
      n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, 
      n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, 
      n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, 
      n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, 
      n15476, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, 
      n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, 
      n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, 
      n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, 
      n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, 
      n15853, n15854, n15855, n15856, n15857, n15858, n15859, n1748, n1747, 
      n1746, n4, n5, n6, n1631, n1633, n1634, n1635, n1636, n1637, n1638, n1639
      , n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, 
      n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, 
      n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, 
      n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, 
      n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, 
      n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
      n1700, n1701, n1703, n1704, n1705, n1707, n1708, n1709, n1711, n1712, 
      n1714, n1715, n1716, n1718, n1719, n1721, n1723, n1725, n1726, n1727, 
      n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, 
      n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1749, n1750, n1751, 
      n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, 
      n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, 
      n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, 
      n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, 
      n1792, n1793, n1794, n1795, n1796, n1797, n1799, n1800, n1801, n1802, 
      n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
      n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
      n1863, n1865, n1867, n1868, n1869, n1870, n1871, n1873, n1874, n1875, 
      n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, 
      n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, 
      n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, 
      n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, 
      n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, 
      n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, 
      n1936, n1937, n1938, n1939, n1940, n1942, n1943, n1945, n1946, n1947, 
      n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, 
      n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, 
      n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, 
      n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, 
      n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, 
      n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, 
      n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2017, n2018, n2019, 
      n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, 
      n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, 
      n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, 
      n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, 
      n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, 
      n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, 
      n2080, n2081, n2082, n2084, n2085, n2086, n2087, n2089, n2090, n2091, 
      n2092, n2093, n2094, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2147, n2150, n2153, n2156, n2159, n2162, n2165, n2168, 
      n2171, n2174, n2177, n2180, n2183, n2186, n2189, n2192, n2198, n2204, 
      n2207, n2213, n2216, n2219, n2222, n2225, n2228, n2231, n2237, n2243, 
      n2249, n2252, n2258, n2261, n2264, n2267, n2270, n2273, n2276, n2279, 
      n2282, n2285, n2288, n2291, n2294, n2297, n2300, n2303, n2306, n2309, 
      n2312, n2315, n2318, n2321, n2324, n2327, n2330, n2333, n2336, n2337, 
      n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, 
      n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, 
      n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, 
      n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2377, n2378, 
      n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, 
      n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, 
      n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, 
      n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, 
      n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, 
      n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, 
      n2439, n2440, n2441, n2443, n2444, n2445, n2446, n2447, n2448, n2449, 
      n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, 
      n2460, n2461, n2462, n2463, n2720, n2721, n2722, n2723, n2724, n2725, 
      n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, 
      n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, 
      n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, 
      n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2766, 
      n2767, n2768, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, 
      n2778, n2779, n2780, n2781, n2782, n2783, n2977, n2979, n2980, n2981, 
      n2982, n2983, n2985, n2986, n2987, n2988, n2990, n2992, n2993, n2994, 
      n2995, n2997, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, 
      n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
      n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, 
      n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
      n3037, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, 
      n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, 
      n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, 
      n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, 
      n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, 
      n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, 
      n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3170, n3172, 
      n3174, n3176, n3178, n3180, n3184, n3186, n3188, n3190, n3192, n3194, 
      n3196, n3198, n3202, n3206, n3208, n3210, n3212, n3214, n3216, n3218, 
      n3220, n3222, n3224, n3226, n3232, n3236, n3242, n3248, n3250, n3252, 
      n3254, n3256, n3258, n3260, n3262, n3264, n3266, n3268, n3270, n3272, 
      n3274, n3276, n3278, n3280, n3282, n3284, n3286, n3288, n3290, n3292, 
      n3294, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3367, n3368, 
      n3369, n3370, n3435, n3436, n3437, n3438, n3503, n3504, n3570, n3571, 
      n3572, n3638, n3639, n3640, n3705, n3706, n3771, n3772, n3837, n3838, 
      n3839, n3906, n3972, n4039, n4106, n4107, n4108, n4109, n4174, n4175, 
      n4176, n4177, n4178, n4243, n4244, n4245, n4310, n4311, n4312, n4377, 
      n4378, n4379, n4380, n4445, n4446, n4447, n4512, n4513, n4514, n4515, 
      n4516, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4652, n4653, 
      n4718, n4719, n4784, n4785, n4786, n4852, n4853, n4854, n4856, n4857, 
      n4922, n4923, n4988, n4989, n5054, n5055, n5056, n5121, n5188, n5254, 
      n5292, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, 
      n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, 
      n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, 
      n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, 
      n5334, n5335, n5337, n5338, n5339, n5341, n5342, n5343, n5344, n5345, 
      n5346, n5347, n5348, n5349, n5350, n5353, n5358, n5362, n5365, n5366, 
      n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, 
      n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, 
      n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, 
      n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5407, 
      n5408, n5409, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, 
      n5419, n5420, n5423, n5427, n5430, n5433, n5434, n5435, n5436, n5437, 
      n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, 
      n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, 
      n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, 
      n5468, n5469, n5470, n5471, n5472, n5473, n5475, n5476, n5477, n5479, 
      n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5493, 
      n5496, n5499, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, 
      n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, 
      n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, 
      n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, 
      n5540, n5541, n5542, n5544, n5545, n5546, n5548, n5549, n5550, n5551, 
      n5552, n5553, n5554, n5555, n5556, n5557, n5563, n5565, n5568, n5571, 
      n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, 
      n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, 
      n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, 
      n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, 
      n5613, n5614, n5615, n5617, n5618, n5619, n5620, n5621, n5622, n5623, 
      n5624, n5625, n5626, n5631, n5633, n5636, n5639, n5640, n5641, n5642, 
      n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, 
      n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, 
      n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, 
      n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5681, n5682, n5683, 
      n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5697, 
      n5701, n5703, n5706, n5709, n5710, n5711, n5712, n5713, n5714, n5715, 
      n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, 
      n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, 
      n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, 
      n5746, n5747, n5748, n5749, n5751, n5752, n5753, n5755, n5756, n5757, 
      n5758, n5759, n5760, n5761, n5762, n5768, n5770, n5773, n5775, n5778, 
      n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, 
      n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, 
      n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, 
      n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, 
      n5821, n5823, n5824, n5825, n5827, n5828, n5829, n5830, n5831, n5832, 
      n5833, n5834, n5836, n5837, n5840, n5842, n5845, n5848, n5849, n5850, 
      n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, 
      n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, 
      n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, 
      n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5890, n5891, 
      n5892, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5902, n5903, 
      n5904, n5907, n5909, n5912, n5915, n5916, n5917, n5918, n5919, n5920, 
      n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, 
      n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, 
      n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, 
      n5951, n5952, n5953, n5954, n5955, n5957, n5958, n5959, n5961, n5962, 
      n5963, n5964, n5965, n5967, n5969, n5970, n5971, n5972, n5975, n5977, 
      n5980, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, 
      n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, 
      n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, 
      n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, 
      n6022, n6023, n6025, n6026, n6027, n6029, n6030, n6031, n6032, n6034, 
      n6036, n6037, n6038, n6039, n6040, n6043, n6045, n6048, n6051, n6052, 
      n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, 
      n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, 
      n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, 
      n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6093, 
      n6094, n6095, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, 
      n6105, n6106, n6109, n6111, n6114, n6117, n6118, n6119, n6120, n6121, 
      n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, 
      n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, 
      n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, 
      n6152, n6153, n6154, n6155, n6156, n6157, n6159, n6160, n6161, n6163, 
      n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6175, 
      n6177, n6180, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, 
      n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, 
      n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, 
      n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, 
      n6221, n6222, n6223, n6225, n6226, n6227, n6229, n6230, n6231, n6232, 
      n6233, n6234, n6235, n6236, n6237, n6238, n6241, n6243, n6246, n6249, 
      n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, 
      n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, 
      n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, 
      n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, 
      n6291, n6292, n6293, n6295, n6296, n6297, n6298, n6299, n6300, n6301, 
      n6302, n6303, n6304, n6307, n6309, n6312, n6315, n6316, n6317, n6318, 
      n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, 
      n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, 
      n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, 
      n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6357, n6358, n6359, 
      n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, 
      n6373, n6375, n6378, n6381, n6382, n6383, n6384, n6385, n6386, n6387, 
      n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, 
      n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, 
      n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, 
      n6418, n6419, n6420, n6421, n6423, n6424, n6425, n6427, n6428, n6429, 
      n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6439, n6441, n6444, 
      n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, 
      n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, 
      n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, 
      n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, 
      n6487, n6489, n6490, n6491, n6493, n6494, n6495, n6496, n6497, n6498, 
      n6499, n6500, n6501, n6502, n6505, n6507, n6510, n6513, n6514, n6515, 
      n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, 
      n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, 
      n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, 
      n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6555, n6556, 
      n6557, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, 
      n6568, n6571, n6573, n6576, n6579, n6580, n6581, n6582, n6583, n6584, 
      n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, 
      n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, 
      n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, 
      n6615, n6616, n6617, n6618, n6619, n6621, n6622, n6623, n6625, n6626, 
      n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6637, n6639, 
      n6642, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, 
      n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, 
      n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, 
      n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, 
      n6685, n6686, n6688, n6689, n6690, n6692, n6693, n6694, n6695, n6697, 
      n6698, n6699, n6700, n6701, n6702, n6705, n6707, n6710, n6713, n6714, 
      n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, 
      n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, 
      n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, 
      n6745, n6746, n6747, n6748, n6750, n6751, n6752, n6753, n6754, n6756, 
      n6757, n6758, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, 
      n6768, n6769, n6772, n6774, n6777, n6780, n6781, n6782, n6783, n6784, 
      n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, 
      n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6803, n6804, n6805, 
      n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, 
      n6816, n6817, n6818, n6819, n6820, n6821, n6823, n6824, n6825, n6827, 
      n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6839, 
      n6841, n6844, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, 
      n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, 
      n6865, n6866, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, 
      n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, 
      n6886, n6887, n6888, n6890, n6891, n6892, n6894, n6895, n6896, n6897, 
      n6898, n6899, n6900, n6901, n6902, n6903, n6906, n6908, n6911, n6914, 
      n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, 
      n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, 
      n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, 
      n6945, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, 
      n6957, n6958, n6959, n6961, n6962, n6963, n6964, n6965, n6966, n6967, 
      n6968, n6969, n6970, n6973, n6975, n6978, n6981, n6982, n6983, n6984, 
      n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, 
      n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, 
      n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, 
      n7015, n7016, n7017, n7018, n7019, n7020, n7021, n9263, n9264, n9266, 
      n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, 
      n9280, n9282, n9285, n9288, n9289, n9290, n9291, n9292, n9293, n9294, 
      n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, 
      n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, 
      n9315, n9316, n9317, n9319, n9320, n9321, n9322, n9323, n9324, n9325, 
      n9326, n9327, n9328, n9329, n9331, n9332, n9333, n9335, n9336, n9337, 
      n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9347, n9349, n9352, 
      n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, 
      n9365, n9366, n9367, n9368, n9369, n9370, n9372, n9373, n9374, n9375, 
      n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, 
      n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, 
      n9396, n9398, n9399, n9400, n9402, n9403, n9404, n9405, n9406, n9407, 
      n9408, n9409, n9410, n9411, n9414, n9416, n9419, n9422, n9423, n9425, 
      n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, 
      n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, 
      n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, 
      n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9465, n9466, 
      n9467, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9478, 
      n9479, n9482, n9484, n9487, n9490, n9491, n9492, n9493, n9494, n9495, 
      n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, 
      n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, 
      n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, 
      n9526, n9527, n9528, n9529, n9531, n9533, n9534, n9535, n9537, n9538, 
      n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9549, n9551, 
      n9554, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, 
      n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, 
      n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9584, n9585, n9586, 
      n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, 
      n9597, n9598, n9600, n9601, n9602, n9604, n9605, n9606, n9607, n9608, 
      n9609, n9610, n9611, n9612, n9613, n9616, n9618, n9621, n9624, n9625, 
      n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, 
      n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, 
      n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, 
      n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9667, 
      n9668, n9669, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, 
      n9679, n9680, n9683, n9685, n9688, n9692, n9693, n9694, n9695, n9696, 
      n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, 
      n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, 
      n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, 
      n9727, n9728, n9729, n9730, n9731, n9732, n9734, n9735, n9736, n9738, 
      n9739, n9740, n9741, n9743, n9744, n9745, n9746, n9747, n9748, n9751, 
      n9753, n9756, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, 
      n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, 
      n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, 
      n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9796, n9797, 
      n9798, n9799, n9800, n9802, n9803, n9804, n9806, n9807, n9808, n9809, 
      n9810, n9811, n9812, n9813, n9814, n9815, n9818, n9820, n9823, n9826, 
      n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, 
      n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, 
      n9847, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, 
      n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, 
      n9869, n9870, n9871, n9873, n9874, n9875, n9876, n9877, n9878, n9879, 
      n9880, n9881, n9882, n9885, n9887, n9890, n9893, n9894, n9895, n9896, 
      n9897, n9898, n9899, n9900, n9902, n9903, n9904, n9905, n9906, n9907, 
      n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, 
      n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, 
      n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9936, n9937, n9938, 
      n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, 
      n9952, n9955, n9958, n9961, n9962, n9963, n9964, n9965, n9966, n9967, 
      n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, 
      n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, 
      n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, 
      n9998, n9999, n10000, n10001, n10003, n10004, n10005, n10008, n10009, 
      n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10020, 
      n10022, n10025, n10028, n10029, n10030, n10031, n10032, n10033, n10034, 
      n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, 
      n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, 
      n10053, n10054, n10055, n10056, n10057, n10058, n10060, n10061, n10062, 
      n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10071, n10072, 
      n10073, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, 
      n10083, n10084, n10087, n10089, n10092, n10095, n10096, n10097, n10098, 
      n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, 
      n10108, n10109, n10110, n10111, n10113, n10114, n10115, n10116, n10117, 
      n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, 
      n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, 
      n10136, n10138, n10139, n10140, n10142, n10143, n10144, n10145, n10146, 
      n10147, n10148, n10149, n10150, n10151, n10154, n10156, n10159, n10162, 
      n10163, n10164, n10166, n10167, n10168, n10169, n10170, n10171, n10172, 
      n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, 
      n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, 
      n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, 
      n10200, n10201, n10202, n10203, n10205, n10206, n10207, n10209, n10210, 
      n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10219, n10222, 
      n10224, n10227, n10230, n10231, n10232, n10233, n10234, n10235, n10236, 
      n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, 
      n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, 
      n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, 
      n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10273, n10274, 
      n10275, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, 
      n10285, n10286, n10289, n10291, n10294, n10297, n10298, n10299, n10300, 
      n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, 
      n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, 
      n10319, n10320, n10321, n10322, n10323, n10325, n10326, n10327, n10328, 
      n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, 
      n10338, n10340, n10341, n10342, n10344, n10345, n10346, n10347, n10348, 
      n10349, n10350, n10351, n10352, n10353, n10356, n10358, n10361, n10364, 
      n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, 
      n10374, n10375, n10376, n10378, n10379, n10380, n10381, n10382, n10383, 
      n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, 
      n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, 
      n10402, n10403, n10404, n10405, n10407, n10408, n10409, n10411, n10412, 
      n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10423, 
      n10425, n10428, n10432, n10433, n10434, n10435, n10436, n10437, n10438, 
      n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, 
      n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, 
      n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, 
      n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10474, n10475, 
      n10476, n10478, n10479, n10480, n10481, n10482, n10484, n10485, n10486, 
      n10487, n10488, n10491, n10493, n10496, n10499, n10500, n10501, n10502, 
      n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, 
      n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, 
      n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, 
      n10530, n10531, n10532, n10533, n10534, n10535, n10537, n10538, n10539, 
      n10540, n10542, n10543, n10544, n10546, n10547, n10548, n10549, n10550, 
      n10551, n10552, n10553, n10554, n10555, n10558, n10560, n10563, n10566, 
      n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, 
      n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, 
      n10585, n10586, n10587, n10588, n10590, n10591, n10592, n10593, n10594, 
      n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, 
      n10604, n10605, n10606, n10607, n10609, n10610, n10611, n10613, n10614, 
      n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10625, 
      n10627, n10630, n10633, n10634, n10635, n10636, n10637, n10638, n10639, 
      n10640, n10641, n10643, n10644, n10645, n10646, n10647, n10648, n10649, 
      n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, 
      n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, 
      n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10676, n10677, 
      n10678, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, 
      n10688, n10689, n10692, n10694, n10698, n10701, n10702, n10703, n10704, 
      n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, 
      n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, 
      n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, 
      n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, 
      n10741, n10743, n10744, n10745, n10747, n10749, n10750, n10751, n10752, 
      n10753, n10754, n10755, n10756, n10757, n10760, n10762, n10765, n10768, 
      n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, 
      n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, 
      n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, 
      n10796, n10797, n10798, n10799, n10800, n10802, n10803, n10804, n10805, 
      n10806, n10807, n10808, n10809, n10811, n10812, n10813, n10815, n10816, 
      n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10827, 
      n10829, n10832, n10835, n10836, n10837, n10838, n10839, n10840, n10841, 
      n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, 
      n10851, n10852, n10853, n10855, n10856, n10857, n10858, n10859, n10860, 
      n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, 
      n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10878, n10879, 
      n10880, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, 
      n10890, n10891, n10894, n10896, n10899, n10902, n10903, n10904, n10905, 
      n10906, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, 
      n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, 
      n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, 
      n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, 
      n10943, n10945, n10946, n10947, n10949, n10950, n10951, n10952, n10953, 
      n10954, n10955, n10956, n10957, n10958, n10962, n10964, n10967, n10970, 
      n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, 
      n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, 
      n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, 
      n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, 
      n11007, n11008, n11009, n11010, n11012, n11014, n11015, n11017, n11018, 
      n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11029, 
      n11031, n11034, n11037, n11038, n11039, n11040, n11041, n11042, n11043, 
      n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, 
      n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, 
      n11062, n11063, n11064, n11065, n11067, n11068, n11069, n11070, n11071, 
      n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11080, n11081, 
      n11082, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, 
      n11092, n11093, n11096, n11098, n11101, n11104, n11105, n11106, n11107, 
      n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, 
      n11117, n11118, n11120, n11121, n11122, n11123, n11124, n11125, n11126, 
      n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, 
      n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, 
      n11145, n11147, n11148, n11149, n11151, n11152, n11153, n11154, n11155, 
      n11156, n11157, n11158, n11159, n11160, n11163, n11165, n11168, n11171, 
      n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, 
      n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, 
      n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, 
      n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, 
      n11209, n11210, n11211, n11212, n11214, n11215, n11216, n11218, n11219, 
      n11220, n11221, n11222, n11223, n11224, n11226, n11227, n11228, n11231, 
      n11233, n11236, n11239, n11240, n11241, n11242, n11243, n11244, n11245, 
      n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, 
      n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, 
      n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, 
      n11273, n11274, n11275, n11276, n11277, n11279, n11280, n11282, n11283, 
      n11284, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, 
      n11294, n11295, n11298, n11300, n11303, n11306, n11307, n11308, n11309, 
      n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, 
      n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, 
      n11328, n11329, n11330, n11332, n11333, n11334, n11335, n11336, n11337, 
      n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, 
      n11347, n11349, n11350, n11351, n11353, n11354, n11355, n11356, n11357, 
      n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, 
      n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, 
      n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11385, 
      n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, 
      n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, 
      n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, 
      n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, 
      n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, 
      n11431, n11432, n11433, n11434, n11435, n11437, n11438, n11439, n11440, 
      n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, 
      n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, 
      n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, 
      n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, 
      n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, 
      n11486, n11487, n11488, n11490, n11491, n11492, n11493, n11494, n11495, 
      n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, 
      n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, 
      n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, 
      n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, 
      n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, 
      n11541, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, 
      n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, 
      n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, 
      n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, 
      n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, 
      n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11596, 
      n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, 
      n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, 
      n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, 
      n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, 
      n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, 
      n11642, n11643, n11644, n11645, n11646, n11647, n11649, n11650, n11651, 
      n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, 
      n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, 
      n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, 
      n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, 
      n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, 
      n11697, n11698, n11699, n11700, n11702, n11703, n11704, n11705, n11706, 
      n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, 
      n11716, n11717, n11718, n11719, n11721, n11722, n11723, n11724, n11725, 
      n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, 
      n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, 
      n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, 
      n11753, n11755, n11756, n11757, n11758, n17696, n17697, n17698, n17699, 
      n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, 
      n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, 
      n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, 
      n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, 
      n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, 
      n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, 
      n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, 
      n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, 
      n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, 
      n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, 
      n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, 
      n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, 
      n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, 
      n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, 
      n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, 
      n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, 
      n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, 
      n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, 
      n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, 
      n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, 
      n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, 
      n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, 
      n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, 
      n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, 
      n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, 
      n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, 
      n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, 
      n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, 
      n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, 
      n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, 
      n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, 
      n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, 
      n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, 
      n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, 
      n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, 
      n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, 
      n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, 
      n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, 
      n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, 
      n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, 
      n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, 
      n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, 
      n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, 
      n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, 
      n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, 
      n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, 
      n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, 
      n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, 
      n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, 
      n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, 
      n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, 
      n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, 
      n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, 
      n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, 
      n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, 
      n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, 
      n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, 
      n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, 
      n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, 
      n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, 
      n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, 
      n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, 
      n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, 
      n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, 
      n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, 
      n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, 
      n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, 
      n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, 
      n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, 
      n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, 
      n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, 
      n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, 
      n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, 
      n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, 
      n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, 
      n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, 
      n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, 
      n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, 
      n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, 
      n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, 
      n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, 
      n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, 
      n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, 
      n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, 
      n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, 
      n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, 
      n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, 
      n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, 
      n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, 
      n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, 
      n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, 
      n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, 
      n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, 
      n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, 
      n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, 
      n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, 
      n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, 
      n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, 
      n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, 
      n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, 
      n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, 
      n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, 
      n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, 
      n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, 
      n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, 
      n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, 
      n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, 
      n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, 
      n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, 
      n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, 
      n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, 
      n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, 
      n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, 
      n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, 
      n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, 
      n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, 
      n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, 
      n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, 
      n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, 
      n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, 
      n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, 
      n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, 
      n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, 
      n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, 
      n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, 
      n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, 
      n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, 
      n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, 
      n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, 
      n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, 
      n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, 
      n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, 
      n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, 
      n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, 
      n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, 
      n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, 
      n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, 
      n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, 
      n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, 
      n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, 
      n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, 
      n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, 
      n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, 
      n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, 
      n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, 
      n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, 
      n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, 
      n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, 
      n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, 
      n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, 
      n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, 
      n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, 
      n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, 
      n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, 
      n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, 
      n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, 
      n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, 
      n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, 
      n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, 
      n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, 
      n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, 
      n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, 
      n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, 
      n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, 
      n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, 
      n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, 
      n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, 
      n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, 
      n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, 
      n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, 
      n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, 
      n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, 
      n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, 
      n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, 
      n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, 
      n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, 
      n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, 
      n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, 
      n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, 
      n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, 
      n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, 
      n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, 
      n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, 
      n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, 
      n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, 
      n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, 
      n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, 
      n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, 
      n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, 
      n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, 
      n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, 
      n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, 
      n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, 
      n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, 
      n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, 
      n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, 
      n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, 
      n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, 
      n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, 
      n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, 
      n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, 
      n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, 
      n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, 
      n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, 
      n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, 
      n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, 
      n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, 
      n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, 
      n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, 
      n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, 
      n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, 
      n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, 
      n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, 
      n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, 
      n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, 
      n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, 
      n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, 
      n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, 
      n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, 
      n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, 
      n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, 
      n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, 
      n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, 
      n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, 
      n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, 
      n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, 
      n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, 
      n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, 
      n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, 
      n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, 
      n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, 
      n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, 
      n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, 
      n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, 
      n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, 
      n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, 
      n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, 
      n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, 
      n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, 
      n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, 
      n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, 
      n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, 
      n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, 
      n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, 
      n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, 
      n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, 
      n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, 
      n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, 
      n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, 
      n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, 
      n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, 
      n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, 
      n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, 
      n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, 
      n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, 
      n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, 
      n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, 
      n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, 
      n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, 
      n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, 
      n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, 
      n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, 
      n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, 
      n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, 
      n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, 
      n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, 
      n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, 
      n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, 
      n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, 
      n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, 
      n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, 
      n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, 
      n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, 
      n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, 
      n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, 
      n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, 
      n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, 
      n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, 
      n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, 
      n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, 
      n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, 
      n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, 
      n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, 
      n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, 
      n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, 
      n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, 
      n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, 
      n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, 
      n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, 
      n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, 
      n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, 
      n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, 
      n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, 
      n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, 
      n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, 
      n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, 
      n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, 
      n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, 
      n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, 
      n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, 
      n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, 
      n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, 
      n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, 
      n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, 
      n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, 
      n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, 
      n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, 
      n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, 
      n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, 
      n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, 
      n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, 
      n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, 
      n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, 
      n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, 
      n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, 
      n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, 
      n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, 
      n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, 
      n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, 
      n20571, n20572, n20573, n20574, n_1006, n_1007, n_1008, n_1009, n_1010, 
      n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, 
      n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125 : std_logic;

begin
   out_to_mem <= ( out_to_mem_63_port, out_to_mem_62_port, out_to_mem_61_port, 
      out_to_mem_60_port, out_to_mem_59_port, out_to_mem_58_port, 
      out_to_mem_57_port, out_to_mem_56_port, out_to_mem_55_port, 
      out_to_mem_54_port, out_to_mem_53_port, out_to_mem_52_port, 
      out_to_mem_51_port, out_to_mem_50_port, out_to_mem_49_port, 
      out_to_mem_48_port, out_to_mem_47_port, out_to_mem_46_port, 
      out_to_mem_45_port, out_to_mem_44_port, out_to_mem_43_port, 
      out_to_mem_42_port, out_to_mem_41_port, out_to_mem_40_port, 
      out_to_mem_39_port, out_to_mem_38_port, out_to_mem_37_port, 
      out_to_mem_36_port, out_to_mem_35_port, out_to_mem_34_port, 
      out_to_mem_33_port, out_to_mem_32_port, out_to_mem_31_port, 
      out_to_mem_30_port, out_to_mem_29_port, out_to_mem_28_port, 
      out_to_mem_27_port, out_to_mem_26_port, out_to_mem_25_port, 
      out_to_mem_24_port, out_to_mem_23_port, out_to_mem_22_port, 
      out_to_mem_21_port, out_to_mem_20_port, out_to_mem_19_port, 
      out_to_mem_18_port, out_to_mem_17_port, out_to_mem_16_port, 
      out_to_mem_15_port, out_to_mem_14_port, out_to_mem_13_port, 
      out_to_mem_12_port, out_to_mem_11_port, out_to_mem_10_port, 
      out_to_mem_9_port, out_to_mem_8_port, out_to_mem_7_port, 
      out_to_mem_6_port, out_to_mem_5_port, out_to_mem_4_port, 
      out_to_mem_3_port, out_to_mem_2_port, out_to_mem_1_port, 
      out_to_mem_0_port );
   
   out2_reg_63_inst : DFF_X1 port map( D => n7277, CK => clk, Q => out2(63), QN
                           => n2335);
   out1_reg_63_inst : DFF_X1 port map( D => n7276, CK => clk, Q => out1(63), QN
                           => n2334);
   out2_reg_62_inst : DFF_X1 port map( D => n7273, CK => clk, Q => out2(62), QN
                           => n2332);
   out1_reg_62_inst : DFF_X1 port map( D => n7272, CK => clk, Q => out1(62), QN
                           => n2331);
   out2_reg_61_inst : DFF_X1 port map( D => n7269, CK => clk, Q => out2(61), QN
                           => n2329);
   out1_reg_61_inst : DFF_X1 port map( D => n7268, CK => clk, Q => out1(61), QN
                           => n2328);
   out2_reg_60_inst : DFF_X1 port map( D => n7265, CK => clk, Q => out2(60), QN
                           => n2326);
   out1_reg_60_inst : DFF_X1 port map( D => n7264, CK => clk, Q => out1(60), QN
                           => n2325);
   out2_reg_59_inst : DFF_X1 port map( D => n7261, CK => clk, Q => out2(59), QN
                           => n2323);
   out1_reg_59_inst : DFF_X1 port map( D => n7260, CK => clk, Q => out1(59), QN
                           => n2322);
   out2_reg_58_inst : DFF_X1 port map( D => n7257, CK => clk, Q => out2(58), QN
                           => n2320);
   out1_reg_58_inst : DFF_X1 port map( D => n7256, CK => clk, Q => out1(58), QN
                           => n2319);
   out2_reg_57_inst : DFF_X1 port map( D => n7253, CK => clk, Q => out2(57), QN
                           => n2317);
   out1_reg_57_inst : DFF_X1 port map( D => n7252, CK => clk, Q => out1(57), QN
                           => n2316);
   out2_reg_56_inst : DFF_X1 port map( D => n7249, CK => clk, Q => out2(56), QN
                           => n2314);
   out1_reg_56_inst : DFF_X1 port map( D => n7248, CK => clk, Q => out1(56), QN
                           => n2313);
   out2_reg_55_inst : DFF_X1 port map( D => n7245, CK => clk, Q => out2(55), QN
                           => n2311);
   out1_reg_55_inst : DFF_X1 port map( D => n7244, CK => clk, Q => out1(55), QN
                           => n2310);
   out2_reg_54_inst : DFF_X1 port map( D => n7241, CK => clk, Q => out2(54), QN
                           => n2308);
   out1_reg_54_inst : DFF_X1 port map( D => n7240, CK => clk, Q => out1(54), QN
                           => n2307);
   out2_reg_53_inst : DFF_X1 port map( D => n7237, CK => clk, Q => out2(53), QN
                           => n2305);
   out1_reg_53_inst : DFF_X1 port map( D => n7236, CK => clk, Q => out1(53), QN
                           => n2304);
   out2_reg_52_inst : DFF_X1 port map( D => n7233, CK => clk, Q => out2(52), QN
                           => n2302);
   out1_reg_52_inst : DFF_X1 port map( D => n7232, CK => clk, Q => out1(52), QN
                           => n2301);
   out2_reg_51_inst : DFF_X1 port map( D => n7229, CK => clk, Q => out2(51), QN
                           => n2299);
   out1_reg_51_inst : DFF_X1 port map( D => n7228, CK => clk, Q => out1(51), QN
                           => n2298);
   out2_reg_50_inst : DFF_X1 port map( D => n7225, CK => clk, Q => out2(50), QN
                           => n2296);
   out1_reg_50_inst : DFF_X1 port map( D => n7224, CK => clk, Q => out1(50), QN
                           => n2295);
   out2_reg_49_inst : DFF_X1 port map( D => n7221, CK => clk, Q => out2(49), QN
                           => n2293);
   out1_reg_49_inst : DFF_X1 port map( D => n7220, CK => clk, Q => out1(49), QN
                           => n2292);
   out2_reg_48_inst : DFF_X1 port map( D => n7217, CK => clk, Q => out2(48), QN
                           => n2290);
   out1_reg_48_inst : DFF_X1 port map( D => n7216, CK => clk, Q => out1(48), QN
                           => n2289);
   out2_reg_47_inst : DFF_X1 port map( D => n7213, CK => clk, Q => out2(47), QN
                           => n2287);
   out1_reg_47_inst : DFF_X1 port map( D => n7212, CK => clk, Q => out1(47), QN
                           => n2286);
   out2_reg_46_inst : DFF_X1 port map( D => n7209, CK => clk, Q => out2(46), QN
                           => n2284);
   out1_reg_46_inst : DFF_X1 port map( D => n7208, CK => clk, Q => out1(46), QN
                           => n2283);
   out2_reg_45_inst : DFF_X1 port map( D => n7205, CK => clk, Q => out2(45), QN
                           => n2281);
   out1_reg_45_inst : DFF_X1 port map( D => n7204, CK => clk, Q => out1(45), QN
                           => n2280);
   out2_reg_44_inst : DFF_X1 port map( D => n7201, CK => clk, Q => out2(44), QN
                           => n2278);
   out1_reg_44_inst : DFF_X1 port map( D => n7200, CK => clk, Q => out1(44), QN
                           => n2277);
   out2_reg_43_inst : DFF_X1 port map( D => n7197, CK => clk, Q => out2(43), QN
                           => n2275);
   out1_reg_43_inst : DFF_X1 port map( D => n7196, CK => clk, Q => out1(43), QN
                           => n2274);
   out2_reg_42_inst : DFF_X1 port map( D => n7193, CK => clk, Q => out2(42), QN
                           => n2272);
   out1_reg_42_inst : DFF_X1 port map( D => n7192, CK => clk, Q => out1(42), QN
                           => n2271);
   out2_reg_41_inst : DFF_X1 port map( D => n7189, CK => clk, Q => out2(41), QN
                           => n2269);
   out1_reg_41_inst : DFF_X1 port map( D => n7188, CK => clk, Q => out1(41), QN
                           => n2268);
   out2_reg_40_inst : DFF_X1 port map( D => n7185, CK => clk, Q => out2(40), QN
                           => n2266);
   out1_reg_40_inst : DFF_X1 port map( D => n7184, CK => clk, Q => out1(40), QN
                           => n2265);
   out2_reg_39_inst : DFF_X1 port map( D => n7181, CK => clk, Q => out2(39), QN
                           => n2263);
   out1_reg_39_inst : DFF_X1 port map( D => n7180, CK => clk, Q => out1(39), QN
                           => n2262);
   out2_reg_38_inst : DFF_X1 port map( D => n7177, CK => clk, Q => out2(38), QN
                           => n2260);
   out1_reg_38_inst : DFF_X1 port map( D => n7176, CK => clk, Q => out1(38), QN
                           => n2259);
   out2_reg_37_inst : DFF_X1 port map( D => n7173, CK => clk, Q => out2(37), QN
                           => n2257);
   out1_reg_37_inst : DFF_X1 port map( D => n7172, CK => clk, Q => out1(37), QN
                           => n2256);
   out2_reg_36_inst : DFF_X1 port map( D => n7169, CK => clk, Q => out2(36), QN
                           => n2254);
   out1_reg_36_inst : DFF_X1 port map( D => n7168, CK => clk, Q => out1(36), QN
                           => n2253);
   out2_reg_35_inst : DFF_X1 port map( D => n7165, CK => clk, Q => out2(35), QN
                           => n2251);
   out1_reg_35_inst : DFF_X1 port map( D => n7164, CK => clk, Q => out1(35), QN
                           => n2250);
   out2_reg_34_inst : DFF_X1 port map( D => n7161, CK => clk, Q => out2(34), QN
                           => n2248);
   out1_reg_34_inst : DFF_X1 port map( D => n7160, CK => clk, Q => out1(34), QN
                           => n2247);
   out2_reg_33_inst : DFF_X1 port map( D => n7157, CK => clk, Q => out2(33), QN
                           => n2245);
   out1_reg_33_inst : DFF_X1 port map( D => n7156, CK => clk, Q => out1(33), QN
                           => n2244);
   out2_reg_32_inst : DFF_X1 port map( D => n7153, CK => clk, Q => out2(32), QN
                           => n2242);
   out1_reg_32_inst : DFF_X1 port map( D => n7152, CK => clk, Q => out1(32), QN
                           => n2241);
   out2_reg_31_inst : DFF_X1 port map( D => n7149, CK => clk, Q => out2(31), QN
                           => n2239);
   out1_reg_31_inst : DFF_X1 port map( D => n7148, CK => clk, Q => out1(31), QN
                           => n2238);
   out2_reg_30_inst : DFF_X1 port map( D => n7145, CK => clk, Q => out2(30), QN
                           => n2236);
   out1_reg_30_inst : DFF_X1 port map( D => n7144, CK => clk, Q => out1(30), QN
                           => n2235);
   out2_reg_29_inst : DFF_X1 port map( D => n7141, CK => clk, Q => out2(29), QN
                           => n2233);
   out1_reg_29_inst : DFF_X1 port map( D => n7140, CK => clk, Q => out1(29), QN
                           => n2232);
   out2_reg_28_inst : DFF_X1 port map( D => n7137, CK => clk, Q => out2(28), QN
                           => n2230);
   out1_reg_28_inst : DFF_X1 port map( D => n7136, CK => clk, Q => out1(28), QN
                           => n2229);
   out2_reg_27_inst : DFF_X1 port map( D => n7133, CK => clk, Q => out2(27), QN
                           => n2227);
   out1_reg_27_inst : DFF_X1 port map( D => n7132, CK => clk, Q => out1(27), QN
                           => n2226);
   out2_reg_26_inst : DFF_X1 port map( D => n7129, CK => clk, Q => out2(26), QN
                           => n2224);
   out1_reg_26_inst : DFF_X1 port map( D => n7128, CK => clk, Q => out1(26), QN
                           => n2223);
   out2_reg_25_inst : DFF_X1 port map( D => n7125, CK => clk, Q => out2(25), QN
                           => n2221);
   out1_reg_25_inst : DFF_X1 port map( D => n7124, CK => clk, Q => out1(25), QN
                           => n2220);
   out2_reg_24_inst : DFF_X1 port map( D => n7121, CK => clk, Q => out2(24), QN
                           => n2218);
   out1_reg_24_inst : DFF_X1 port map( D => n7120, CK => clk, Q => out1(24), QN
                           => n2217);
   out2_reg_23_inst : DFF_X1 port map( D => n7117, CK => clk, Q => out2(23), QN
                           => n2215);
   out1_reg_23_inst : DFF_X1 port map( D => n7116, CK => clk, Q => out1(23), QN
                           => n2214);
   out2_reg_22_inst : DFF_X1 port map( D => n7113, CK => clk, Q => out2(22), QN
                           => n2212);
   out1_reg_22_inst : DFF_X1 port map( D => n7112, CK => clk, Q => out1(22), QN
                           => n2211);
   out2_reg_21_inst : DFF_X1 port map( D => n7109, CK => clk, Q => out2(21), QN
                           => n2209);
   out1_reg_21_inst : DFF_X1 port map( D => n7108, CK => clk, Q => out1(21), QN
                           => n2208);
   out2_reg_20_inst : DFF_X1 port map( D => n7105, CK => clk, Q => out2(20), QN
                           => n2206);
   out1_reg_20_inst : DFF_X1 port map( D => n7104, CK => clk, Q => out1(20), QN
                           => n2205);
   out2_reg_19_inst : DFF_X1 port map( D => n7101, CK => clk, Q => out2(19), QN
                           => n2203);
   out1_reg_19_inst : DFF_X1 port map( D => n7100, CK => clk, Q => out1(19), QN
                           => n2202);
   out2_reg_18_inst : DFF_X1 port map( D => n7097, CK => clk, Q => out2(18), QN
                           => n2200);
   out1_reg_18_inst : DFF_X1 port map( D => n7096, CK => clk, Q => out1(18), QN
                           => n2199);
   out2_reg_17_inst : DFF_X1 port map( D => n7093, CK => clk, Q => out2(17), QN
                           => n2197);
   out1_reg_17_inst : DFF_X1 port map( D => n7092, CK => clk, Q => out1(17), QN
                           => n2196);
   out2_reg_16_inst : DFF_X1 port map( D => n7089, CK => clk, Q => out2(16), QN
                           => n2194);
   out1_reg_16_inst : DFF_X1 port map( D => n7088, CK => clk, Q => out1(16), QN
                           => n2193);
   out2_reg_15_inst : DFF_X1 port map( D => n7085, CK => clk, Q => out2(15), QN
                           => n2191);
   out1_reg_15_inst : DFF_X1 port map( D => n7084, CK => clk, Q => out1(15), QN
                           => n2190);
   out2_reg_14_inst : DFF_X1 port map( D => n7081, CK => clk, Q => out2(14), QN
                           => n2188);
   out1_reg_14_inst : DFF_X1 port map( D => n7080, CK => clk, Q => out1(14), QN
                           => n2187);
   out2_reg_13_inst : DFF_X1 port map( D => n7077, CK => clk, Q => out2(13), QN
                           => n2185);
   out1_reg_13_inst : DFF_X1 port map( D => n7076, CK => clk, Q => out1(13), QN
                           => n2184);
   out2_reg_12_inst : DFF_X1 port map( D => n7073, CK => clk, Q => out2(12), QN
                           => n2182);
   out1_reg_12_inst : DFF_X1 port map( D => n7072, CK => clk, Q => out1(12), QN
                           => n2181);
   out2_reg_11_inst : DFF_X1 port map( D => n7069, CK => clk, Q => out2(11), QN
                           => n2179);
   out1_reg_11_inst : DFF_X1 port map( D => n7068, CK => clk, Q => out1(11), QN
                           => n2178);
   out2_reg_10_inst : DFF_X1 port map( D => n7065, CK => clk, Q => out2(10), QN
                           => n2176);
   out1_reg_10_inst : DFF_X1 port map( D => n7064, CK => clk, Q => out1(10), QN
                           => n2175);
   out2_reg_9_inst : DFF_X1 port map( D => n7061, CK => clk, Q => out2(9), QN 
                           => n2173);
   out1_reg_9_inst : DFF_X1 port map( D => n7060, CK => clk, Q => out1(9), QN 
                           => n2172);
   out2_reg_8_inst : DFF_X1 port map( D => n7057, CK => clk, Q => out2(8), QN 
                           => n2170);
   out1_reg_8_inst : DFF_X1 port map( D => n7056, CK => clk, Q => out1(8), QN 
                           => n2169);
   out2_reg_7_inst : DFF_X1 port map( D => n7053, CK => clk, Q => out2(7), QN 
                           => n2167);
   out1_reg_7_inst : DFF_X1 port map( D => n7052, CK => clk, Q => out1(7), QN 
                           => n2166);
   out2_reg_6_inst : DFF_X1 port map( D => n7049, CK => clk, Q => out2(6), QN 
                           => n2164);
   out1_reg_6_inst : DFF_X1 port map( D => n7048, CK => clk, Q => out1(6), QN 
                           => n2163);
   out2_reg_5_inst : DFF_X1 port map( D => n7045, CK => clk, Q => out2(5), QN 
                           => n2161);
   out1_reg_5_inst : DFF_X1 port map( D => n7044, CK => clk, Q => out1(5), QN 
                           => n2160);
   out2_reg_4_inst : DFF_X1 port map( D => n7041, CK => clk, Q => out2(4), QN 
                           => n2158);
   out1_reg_4_inst : DFF_X1 port map( D => n7040, CK => clk, Q => out1(4), QN 
                           => n2157);
   out2_reg_3_inst : DFF_X1 port map( D => n7037, CK => clk, Q => out2(3), QN 
                           => n2155);
   out1_reg_3_inst : DFF_X1 port map( D => n7036, CK => clk, Q => out1(3), QN 
                           => n2154);
   out2_reg_2_inst : DFF_X1 port map( D => n7033, CK => clk, Q => out2(2), QN 
                           => n2152);
   out1_reg_2_inst : DFF_X1 port map( D => n7032, CK => clk, Q => out1(2), QN 
                           => n2151);
   out2_reg_1_inst : DFF_X1 port map( D => n7029, CK => clk, Q => out2(1), QN 
                           => n2149);
   out1_reg_1_inst : DFF_X1 port map( D => n7028, CK => clk, Q => out1(1), QN 
                           => n2148);
   out2_reg_0_inst : DFF_X1 port map( D => n7025, CK => clk, Q => out2(0), QN 
                           => n2146);
   out1_reg_0_inst : DFF_X1 port map( D => n7024, CK => clk, Q => out1(0), QN 
                           => n2145);
   registers_reg_26_63_inst : DFF_X1 port map( D => n8942, CK => clk, Q => 
                           n_1006, QN => n3574);
   registers_reg_26_62_inst : DFF_X1 port map( D => n8941, CK => clk, Q => 
                           n_1007, QN => n3575);
   registers_reg_26_61_inst : DFF_X1 port map( D => n8940, CK => clk, Q => 
                           n_1008, QN => n3576);
   registers_reg_26_60_inst : DFF_X1 port map( D => n8939, CK => clk, Q => 
                           n_1009, QN => n3577);
   registers_reg_26_59_inst : DFF_X1 port map( D => n8938, CK => clk, Q => 
                           n_1010, QN => n3578);
   registers_reg_26_58_inst : DFF_X1 port map( D => n8937, CK => clk, Q => 
                           n_1011, QN => n3579);
   registers_reg_26_57_inst : DFF_X1 port map( D => n8936, CK => clk, Q => 
                           n_1012, QN => n3580);
   registers_reg_26_56_inst : DFF_X1 port map( D => n8935, CK => clk, Q => 
                           n_1013, QN => n3581);
   registers_reg_26_55_inst : DFF_X1 port map( D => n8934, CK => clk, Q => 
                           n_1014, QN => n3582);
   registers_reg_26_54_inst : DFF_X1 port map( D => n8933, CK => clk, Q => 
                           n_1015, QN => n3583);
   registers_reg_26_53_inst : DFF_X1 port map( D => n8932, CK => clk, Q => 
                           n_1016, QN => n3584);
   registers_reg_26_52_inst : DFF_X1 port map( D => n8931, CK => clk, Q => 
                           n_1017, QN => n3585);
   registers_reg_26_51_inst : DFF_X1 port map( D => n8930, CK => clk, Q => 
                           n_1018, QN => n3586);
   registers_reg_26_50_inst : DFF_X1 port map( D => n8929, CK => clk, Q => 
                           n_1019, QN => n3587);
   registers_reg_26_49_inst : DFF_X1 port map( D => n8928, CK => clk, Q => 
                           n_1020, QN => n3588);
   registers_reg_26_48_inst : DFF_X1 port map( D => n8927, CK => clk, Q => 
                           n_1021, QN => n3589);
   registers_reg_26_47_inst : DFF_X1 port map( D => n8926, CK => clk, Q => 
                           n_1022, QN => n3590);
   registers_reg_26_46_inst : DFF_X1 port map( D => n8925, CK => clk, Q => 
                           n_1023, QN => n3591);
   registers_reg_26_45_inst : DFF_X1 port map( D => n8924, CK => clk, Q => 
                           n_1024, QN => n3592);
   registers_reg_26_44_inst : DFF_X1 port map( D => n8923, CK => clk, Q => 
                           n_1025, QN => n3593);
   registers_reg_26_43_inst : DFF_X1 port map( D => n8922, CK => clk, Q => 
                           n_1026, QN => n3594);
   registers_reg_26_42_inst : DFF_X1 port map( D => n8921, CK => clk, Q => 
                           n_1027, QN => n3595);
   registers_reg_26_41_inst : DFF_X1 port map( D => n8920, CK => clk, Q => 
                           n_1028, QN => n3596);
   registers_reg_26_40_inst : DFF_X1 port map( D => n8919, CK => clk, Q => 
                           n_1029, QN => n3597);
   registers_reg_26_39_inst : DFF_X1 port map( D => n8918, CK => clk, Q => 
                           n_1030, QN => n3598);
   registers_reg_26_38_inst : DFF_X1 port map( D => n8917, CK => clk, Q => 
                           n_1031, QN => n3599);
   registers_reg_26_37_inst : DFF_X1 port map( D => n8916, CK => clk, Q => 
                           n_1032, QN => n3600);
   registers_reg_26_36_inst : DFF_X1 port map( D => n8915, CK => clk, Q => 
                           n_1033, QN => n3601);
   registers_reg_26_35_inst : DFF_X1 port map( D => n8914, CK => clk, Q => 
                           n_1034, QN => n3602);
   registers_reg_26_34_inst : DFF_X1 port map( D => n8913, CK => clk, Q => 
                           n_1035, QN => n3603);
   registers_reg_26_33_inst : DFF_X1 port map( D => n8912, CK => clk, Q => 
                           n_1036, QN => n3604);
   registers_reg_26_32_inst : DFF_X1 port map( D => n8911, CK => clk, Q => 
                           n_1037, QN => n3605);
   registers_reg_26_31_inst : DFF_X1 port map( D => n8910, CK => clk, Q => 
                           n_1038, QN => n3606);
   registers_reg_26_30_inst : DFF_X1 port map( D => n8909, CK => clk, Q => 
                           n_1039, QN => n3607);
   registers_reg_26_29_inst : DFF_X1 port map( D => n8908, CK => clk, Q => 
                           n_1040, QN => n3608);
   registers_reg_26_28_inst : DFF_X1 port map( D => n8907, CK => clk, Q => 
                           n_1041, QN => n3609);
   registers_reg_26_27_inst : DFF_X1 port map( D => n8906, CK => clk, Q => 
                           n_1042, QN => n3610);
   registers_reg_26_26_inst : DFF_X1 port map( D => n8905, CK => clk, Q => 
                           n_1043, QN => n3611);
   registers_reg_26_25_inst : DFF_X1 port map( D => n8904, CK => clk, Q => 
                           n_1044, QN => n3612);
   registers_reg_26_24_inst : DFF_X1 port map( D => n8903, CK => clk, Q => 
                           n_1045, QN => n3613);
   registers_reg_26_23_inst : DFF_X1 port map( D => n8902, CK => clk, Q => 
                           n_1046, QN => n3614);
   registers_reg_26_22_inst : DFF_X1 port map( D => n8901, CK => clk, Q => 
                           n_1047, QN => n3615);
   registers_reg_26_21_inst : DFF_X1 port map( D => n8900, CK => clk, Q => 
                           n_1048, QN => n3616);
   registers_reg_26_20_inst : DFF_X1 port map( D => n8899, CK => clk, Q => 
                           n_1049, QN => n3617);
   registers_reg_26_19_inst : DFF_X1 port map( D => n8898, CK => clk, Q => 
                           n_1050, QN => n3618);
   registers_reg_26_18_inst : DFF_X1 port map( D => n8897, CK => clk, Q => 
                           n_1051, QN => n3619);
   registers_reg_26_17_inst : DFF_X1 port map( D => n8896, CK => clk, Q => 
                           n_1052, QN => n3620);
   registers_reg_26_16_inst : DFF_X1 port map( D => n8895, CK => clk, Q => 
                           n_1053, QN => n3621);
   registers_reg_26_15_inst : DFF_X1 port map( D => n8894, CK => clk, Q => 
                           n_1054, QN => n3622);
   registers_reg_26_14_inst : DFF_X1 port map( D => n8893, CK => clk, Q => 
                           n_1055, QN => n3623);
   registers_reg_26_13_inst : DFF_X1 port map( D => n8892, CK => clk, Q => 
                           n_1056, QN => n3624);
   registers_reg_26_12_inst : DFF_X1 port map( D => n8891, CK => clk, Q => 
                           n_1057, QN => n3625);
   registers_reg_26_11_inst : DFF_X1 port map( D => n8890, CK => clk, Q => 
                           n_1058, QN => n3626);
   registers_reg_26_10_inst : DFF_X1 port map( D => n8889, CK => clk, Q => 
                           n_1059, QN => n3627);
   registers_reg_26_9_inst : DFF_X1 port map( D => n8888, CK => clk, Q => 
                           n_1060, QN => n3628);
   registers_reg_26_8_inst : DFF_X1 port map( D => n8887, CK => clk, Q => 
                           n_1061, QN => n3629);
   registers_reg_26_7_inst : DFF_X1 port map( D => n8886, CK => clk, Q => 
                           n_1062, QN => n3630);
   registers_reg_26_6_inst : DFF_X1 port map( D => n8885, CK => clk, Q => 
                           n_1063, QN => n3631);
   registers_reg_26_5_inst : DFF_X1 port map( D => n8884, CK => clk, Q => 
                           n_1064, QN => n3632);
   registers_reg_26_4_inst : DFF_X1 port map( D => n8883, CK => clk, Q => 
                           n_1065, QN => n3633);
   registers_reg_27_63_inst : DFF_X1 port map( D => n9006, CK => clk, Q => 
                           n18120, QN => n3506);
   registers_reg_27_62_inst : DFF_X1 port map( D => n9005, CK => clk, Q => 
                           n18119, QN => n3507);
   registers_reg_27_61_inst : DFF_X1 port map( D => n9004, CK => clk, Q => 
                           n18118, QN => n3508);
   registers_reg_27_60_inst : DFF_X1 port map( D => n9003, CK => clk, Q => 
                           n18117, QN => n3509);
   registers_reg_27_59_inst : DFF_X1 port map( D => n9002, CK => clk, Q => 
                           n18141, QN => n3510);
   registers_reg_27_58_inst : DFF_X1 port map( D => n9001, CK => clk, Q => 
                           n18140, QN => n3511);
   registers_reg_27_57_inst : DFF_X1 port map( D => n9000, CK => clk, Q => 
                           n18139, QN => n3512);
   registers_reg_27_56_inst : DFF_X1 port map( D => n8999, CK => clk, Q => 
                           n18138, QN => n3513);
   registers_reg_27_55_inst : DFF_X1 port map( D => n8998, CK => clk, Q => 
                           n18137, QN => n3514);
   registers_reg_27_54_inst : DFF_X1 port map( D => n8997, CK => clk, Q => 
                           n18136, QN => n3515);
   registers_reg_27_53_inst : DFF_X1 port map( D => n8996, CK => clk, Q => 
                           n18135, QN => n3516);
   registers_reg_27_52_inst : DFF_X1 port map( D => n8995, CK => clk, Q => 
                           n18134, QN => n3517);
   registers_reg_27_51_inst : DFF_X1 port map( D => n8994, CK => clk, Q => 
                           n18133, QN => n3518);
   registers_reg_27_50_inst : DFF_X1 port map( D => n8993, CK => clk, Q => 
                           n18132, QN => n3519);
   registers_reg_27_49_inst : DFF_X1 port map( D => n8992, CK => clk, Q => 
                           n18131, QN => n3520);
   registers_reg_27_48_inst : DFF_X1 port map( D => n8991, CK => clk, Q => 
                           n18130, QN => n3521);
   registers_reg_27_47_inst : DFF_X1 port map( D => n8990, CK => clk, Q => 
                           n18129, QN => n3522);
   registers_reg_27_46_inst : DFF_X1 port map( D => n8989, CK => clk, Q => 
                           n18128, QN => n3523);
   registers_reg_27_45_inst : DFF_X1 port map( D => n8988, CK => clk, Q => 
                           n18127, QN => n3524);
   registers_reg_27_44_inst : DFF_X1 port map( D => n8987, CK => clk, Q => 
                           n18126, QN => n3525);
   registers_reg_27_43_inst : DFF_X1 port map( D => n8986, CK => clk, Q => 
                           n18125, QN => n3526);
   registers_reg_27_42_inst : DFF_X1 port map( D => n8985, CK => clk, Q => 
                           n18124, QN => n3527);
   registers_reg_27_41_inst : DFF_X1 port map( D => n8984, CK => clk, Q => 
                           n18123, QN => n3528);
   registers_reg_27_40_inst : DFF_X1 port map( D => n8983, CK => clk, Q => 
                           n18122, QN => n3529);
   registers_reg_27_39_inst : DFF_X1 port map( D => n8982, CK => clk, Q => 
                           n18121, QN => n3530);
   registers_reg_27_38_inst : DFF_X1 port map( D => n8981, CK => clk, Q => 
                           n18116, QN => n3531);
   registers_reg_27_37_inst : DFF_X1 port map( D => n8980, CK => clk, Q => 
                           n18175, QN => n3532);
   registers_reg_27_36_inst : DFF_X1 port map( D => n8979, CK => clk, Q => 
                           n18174, QN => n3533);
   registers_reg_27_35_inst : DFF_X1 port map( D => n8978, CK => clk, Q => 
                           n18173, QN => n3534);
   registers_reg_27_34_inst : DFF_X1 port map( D => n8977, CK => clk, Q => 
                           n18172, QN => n3535);
   registers_reg_27_33_inst : DFF_X1 port map( D => n8976, CK => clk, Q => 
                           n18171, QN => n3536);
   registers_reg_27_32_inst : DFF_X1 port map( D => n8975, CK => clk, Q => 
                           n18170, QN => n3537);
   registers_reg_27_31_inst : DFF_X1 port map( D => n8974, CK => clk, Q => 
                           n18169, QN => n3538);
   registers_reg_27_30_inst : DFF_X1 port map( D => n8973, CK => clk, Q => 
                           n18168, QN => n3539);
   registers_reg_27_29_inst : DFF_X1 port map( D => n8972, CK => clk, Q => 
                           n18167, QN => n3540);
   registers_reg_27_28_inst : DFF_X1 port map( D => n8971, CK => clk, Q => 
                           n18166, QN => n3541);
   registers_reg_27_27_inst : DFF_X1 port map( D => n8970, CK => clk, Q => 
                           n18165, QN => n3542);
   registers_reg_27_26_inst : DFF_X1 port map( D => n8969, CK => clk, Q => 
                           n18164, QN => n3543);
   registers_reg_27_25_inst : DFF_X1 port map( D => n8968, CK => clk, Q => 
                           n18163, QN => n3544);
   registers_reg_27_24_inst : DFF_X1 port map( D => n8967, CK => clk, Q => 
                           n18162, QN => n3545);
   registers_reg_27_23_inst : DFF_X1 port map( D => n8966, CK => clk, Q => 
                           n18161, QN => n3546);
   registers_reg_27_22_inst : DFF_X1 port map( D => n8965, CK => clk, Q => 
                           n18160, QN => n3547);
   registers_reg_27_21_inst : DFF_X1 port map( D => n8964, CK => clk, Q => 
                           n18159, QN => n3548);
   registers_reg_27_20_inst : DFF_X1 port map( D => n8963, CK => clk, Q => 
                           n18158, QN => n3549);
   registers_reg_27_19_inst : DFF_X1 port map( D => n8962, CK => clk, Q => 
                           n18157, QN => n3550);
   registers_reg_27_18_inst : DFF_X1 port map( D => n8961, CK => clk, Q => 
                           n18156, QN => n3551);
   registers_reg_27_17_inst : DFF_X1 port map( D => n8960, CK => clk, Q => 
                           n18155, QN => n3552);
   registers_reg_27_16_inst : DFF_X1 port map( D => n8959, CK => clk, Q => 
                           n18154, QN => n3553);
   registers_reg_27_15_inst : DFF_X1 port map( D => n8958, CK => clk, Q => 
                           n18153, QN => n3554);
   registers_reg_27_14_inst : DFF_X1 port map( D => n8957, CK => clk, Q => 
                           n18152, QN => n3555);
   registers_reg_27_13_inst : DFF_X1 port map( D => n8956, CK => clk, Q => 
                           n18151, QN => n3556);
   registers_reg_27_12_inst : DFF_X1 port map( D => n8955, CK => clk, Q => 
                           n18150, QN => n3557);
   registers_reg_27_11_inst : DFF_X1 port map( D => n8954, CK => clk, Q => 
                           n18149, QN => n3558);
   registers_reg_27_10_inst : DFF_X1 port map( D => n8953, CK => clk, Q => 
                           n18148, QN => n3559);
   registers_reg_27_9_inst : DFF_X1 port map( D => n8952, CK => clk, Q => 
                           n18147, QN => n3560);
   registers_reg_27_8_inst : DFF_X1 port map( D => n8951, CK => clk, Q => 
                           n18146, QN => n3561);
   registers_reg_27_7_inst : DFF_X1 port map( D => n8950, CK => clk, Q => 
                           n18145, QN => n3562);
   registers_reg_27_6_inst : DFF_X1 port map( D => n8949, CK => clk, Q => 
                           n18144, QN => n3563);
   registers_reg_27_5_inst : DFF_X1 port map( D => n8948, CK => clk, Q => 
                           n18143, QN => n3564);
   registers_reg_27_4_inst : DFF_X1 port map( D => n8947, CK => clk, Q => 
                           n18142, QN => n3565);
   registers_reg_31_63_inst : DFF_X1 port map( D => n9262, CK => clk, Q => 
                           n18107, QN => n3169);
   registers_reg_31_62_inst : DFF_X1 port map( D => n9261, CK => clk, Q => 
                           n18106, QN => n3171);
   registers_reg_31_61_inst : DFF_X1 port map( D => n9260, CK => clk, Q => 
                           n18105, QN => n3173);
   registers_reg_31_60_inst : DFF_X1 port map( D => n9259, CK => clk, Q => 
                           n18104, QN => n3175);
   registers_reg_31_59_inst : DFF_X1 port map( D => n9258, CK => clk, Q => 
                           n18103, QN => n3177);
   registers_reg_31_58_inst : DFF_X1 port map( D => n9257, CK => clk, Q => 
                           n18102, QN => n3179);
   registers_reg_31_57_inst : DFF_X1 port map( D => n9256, CK => clk, Q => 
                           n18101, QN => n3181);
   registers_reg_31_56_inst : DFF_X1 port map( D => n9255, CK => clk, Q => 
                           n18100, QN => n3183);
   registers_reg_31_55_inst : DFF_X1 port map( D => n9254, CK => clk, Q => 
                           n18099, QN => n3185);
   registers_reg_31_54_inst : DFF_X1 port map( D => n9253, CK => clk, Q => 
                           n18098, QN => n3187);
   registers_reg_31_53_inst : DFF_X1 port map( D => n9252, CK => clk, Q => 
                           n18097, QN => n3189);
   registers_reg_31_52_inst : DFF_X1 port map( D => n9251, CK => clk, Q => 
                           n18096, QN => n3191);
   registers_reg_31_51_inst : DFF_X1 port map( D => n9250, CK => clk, Q => 
                           n18095, QN => n3193);
   registers_reg_31_50_inst : DFF_X1 port map( D => n9249, CK => clk, Q => 
                           n18094, QN => n3195);
   registers_reg_31_49_inst : DFF_X1 port map( D => n9248, CK => clk, Q => 
                           n18093, QN => n3197);
   registers_reg_31_48_inst : DFF_X1 port map( D => n9247, CK => clk, Q => 
                           n18092, QN => n3199);
   registers_reg_31_47_inst : DFF_X1 port map( D => n9246, CK => clk, Q => 
                           n18091, QN => n3201);
   registers_reg_31_46_inst : DFF_X1 port map( D => n9245, CK => clk, Q => 
                           n18090, QN => n3203);
   registers_reg_31_45_inst : DFF_X1 port map( D => n9244, CK => clk, Q => 
                           n18089, QN => n3205);
   registers_reg_31_44_inst : DFF_X1 port map( D => n9243, CK => clk, Q => 
                           n18088, QN => n3207);
   registers_reg_31_43_inst : DFF_X1 port map( D => n9242, CK => clk, Q => 
                           n18087, QN => n3209);
   registers_reg_31_42_inst : DFF_X1 port map( D => n9241, CK => clk, Q => 
                           n18086, QN => n3211);
   registers_reg_31_41_inst : DFF_X1 port map( D => n9240, CK => clk, Q => 
                           n18085, QN => n3213);
   registers_reg_31_40_inst : DFF_X1 port map( D => n9239, CK => clk, Q => 
                           n18084, QN => n3215);
   registers_reg_31_39_inst : DFF_X1 port map( D => n9238, CK => clk, Q => 
                           n18083, QN => n3217);
   registers_reg_31_38_inst : DFF_X1 port map( D => n9237, CK => clk, Q => 
                           n18082, QN => n3219);
   registers_reg_31_37_inst : DFF_X1 port map( D => n9236, CK => clk, Q => 
                           n18081, QN => n3221);
   registers_reg_31_36_inst : DFF_X1 port map( D => n9235, CK => clk, Q => 
                           n18080, QN => n3223);
   registers_reg_31_35_inst : DFF_X1 port map( D => n9234, CK => clk, Q => 
                           n18079, QN => n3225);
   registers_reg_31_34_inst : DFF_X1 port map( D => n9233, CK => clk, Q => 
                           n18078, QN => n3227);
   registers_reg_31_33_inst : DFF_X1 port map( D => n9232, CK => clk, Q => 
                           n18077, QN => n3229);
   registers_reg_31_32_inst : DFF_X1 port map( D => n9231, CK => clk, Q => 
                           n18076, QN => n3231);
   registers_reg_31_31_inst : DFF_X1 port map( D => n9230, CK => clk, Q => 
                           n18075, QN => n3233);
   registers_reg_31_30_inst : DFF_X1 port map( D => n9229, CK => clk, Q => 
                           n18074, QN => n3235);
   registers_reg_31_29_inst : DFF_X1 port map( D => n9228, CK => clk, Q => 
                           n18073, QN => n3237);
   registers_reg_31_28_inst : DFF_X1 port map( D => n9227, CK => clk, Q => 
                           n18072, QN => n3239);
   registers_reg_31_27_inst : DFF_X1 port map( D => n9226, CK => clk, Q => 
                           n18071, QN => n3241);
   registers_reg_31_26_inst : DFF_X1 port map( D => n9225, CK => clk, Q => 
                           n18070, QN => n3243);
   registers_reg_31_25_inst : DFF_X1 port map( D => n9224, CK => clk, Q => 
                           n18069, QN => n3245);
   registers_reg_31_24_inst : DFF_X1 port map( D => n9223, CK => clk, Q => 
                           n18068, QN => n3247);
   registers_reg_31_23_inst : DFF_X1 port map( D => n9222, CK => clk, Q => 
                           n18067, QN => n3249);
   registers_reg_31_22_inst : DFF_X1 port map( D => n9221, CK => clk, Q => 
                           n18066, QN => n3251);
   registers_reg_31_21_inst : DFF_X1 port map( D => n9220, CK => clk, Q => 
                           n18065, QN => n3253);
   registers_reg_31_20_inst : DFF_X1 port map( D => n9219, CK => clk, Q => 
                           n18064, QN => n3255);
   registers_reg_31_19_inst : DFF_X1 port map( D => n9218, CK => clk, Q => 
                           n18063, QN => n3257);
   registers_reg_31_18_inst : DFF_X1 port map( D => n9217, CK => clk, Q => 
                           n18062, QN => n3259);
   registers_reg_31_17_inst : DFF_X1 port map( D => n9216, CK => clk, Q => 
                           n18061, QN => n3261);
   registers_reg_31_16_inst : DFF_X1 port map( D => n9215, CK => clk, Q => 
                           n18060, QN => n3263);
   registers_reg_31_15_inst : DFF_X1 port map( D => n9214, CK => clk, Q => 
                           n18059, QN => n3265);
   registers_reg_31_14_inst : DFF_X1 port map( D => n9213, CK => clk, Q => 
                           n18058, QN => n3267);
   registers_reg_31_13_inst : DFF_X1 port map( D => n9212, CK => clk, Q => 
                           n18057, QN => n3269);
   registers_reg_31_12_inst : DFF_X1 port map( D => n9211, CK => clk, Q => 
                           n18056, QN => n3271);
   registers_reg_31_11_inst : DFF_X1 port map( D => n9210, CK => clk, Q => 
                           n18115, QN => n3273);
   registers_reg_31_10_inst : DFF_X1 port map( D => n9209, CK => clk, Q => 
                           n18114, QN => n3275);
   registers_reg_31_9_inst : DFF_X1 port map( D => n9208, CK => clk, Q => 
                           n18113, QN => n3277);
   registers_reg_31_8_inst : DFF_X1 port map( D => n9207, CK => clk, Q => 
                           n18112, QN => n3279);
   registers_reg_31_7_inst : DFF_X1 port map( D => n9206, CK => clk, Q => 
                           n18111, QN => n3281);
   registers_reg_31_6_inst : DFF_X1 port map( D => n9205, CK => clk, Q => 
                           n18110, QN => n3283);
   registers_reg_31_5_inst : DFF_X1 port map( D => n9204, CK => clk, Q => 
                           n18109, QN => n3285);
   registers_reg_31_4_inst : DFF_X1 port map( D => n9203, CK => clk, Q => 
                           n18108, QN => n3287);
   registers_reg_19_63_inst : DFF_X1 port map( D => n8494, CK => clk, Q => 
                           n17795, QN => n4040);
   registers_reg_19_62_inst : DFF_X1 port map( D => n8493, CK => clk, Q => 
                           n17794, QN => n4041);
   registers_reg_19_61_inst : DFF_X1 port map( D => n8492, CK => clk, Q => 
                           n17793, QN => n4042);
   registers_reg_19_60_inst : DFF_X1 port map( D => n8491, CK => clk, Q => 
                           n17792, QN => n4043);
   registers_reg_19_59_inst : DFF_X1 port map( D => n8490, CK => clk, Q => 
                           n17767, QN => n4044);
   registers_reg_19_58_inst : DFF_X1 port map( D => n8489, CK => clk, Q => 
                           n17766, QN => n4045);
   registers_reg_19_57_inst : DFF_X1 port map( D => n8488, CK => clk, Q => 
                           n17765, QN => n4046);
   registers_reg_19_56_inst : DFF_X1 port map( D => n8487, CK => clk, Q => 
                           n17764, QN => n4047);
   registers_reg_19_55_inst : DFF_X1 port map( D => n8486, CK => clk, Q => 
                           n17763, QN => n4048);
   registers_reg_19_54_inst : DFF_X1 port map( D => n8485, CK => clk, Q => 
                           n17762, QN => n4049);
   registers_reg_19_53_inst : DFF_X1 port map( D => n8484, CK => clk, Q => 
                           n17761, QN => n4050);
   registers_reg_19_52_inst : DFF_X1 port map( D => n8483, CK => clk, Q => 
                           n17760, QN => n4051);
   registers_reg_19_51_inst : DFF_X1 port map( D => n8482, CK => clk, Q => 
                           n17759, QN => n4052);
   registers_reg_19_50_inst : DFF_X1 port map( D => n8481, CK => clk, Q => 
                           n17758, QN => n4053);
   registers_reg_19_49_inst : DFF_X1 port map( D => n8480, CK => clk, Q => 
                           n17757, QN => n4054);
   registers_reg_19_48_inst : DFF_X1 port map( D => n8479, CK => clk, Q => 
                           n17756, QN => n4055);
   registers_reg_19_47_inst : DFF_X1 port map( D => n8478, CK => clk, Q => 
                           n17804, QN => n4056);
   registers_reg_19_46_inst : DFF_X1 port map( D => n8477, CK => clk, Q => 
                           n17803, QN => n4057);
   registers_reg_19_45_inst : DFF_X1 port map( D => n8476, CK => clk, Q => 
                           n17802, QN => n4058);
   registers_reg_19_44_inst : DFF_X1 port map( D => n8475, CK => clk, Q => 
                           n17801, QN => n4059);
   registers_reg_19_43_inst : DFF_X1 port map( D => n8474, CK => clk, Q => 
                           n17800, QN => n4060);
   registers_reg_19_42_inst : DFF_X1 port map( D => n8473, CK => clk, Q => 
                           n17799, QN => n4061);
   registers_reg_19_41_inst : DFF_X1 port map( D => n8472, CK => clk, Q => 
                           n17798, QN => n4062);
   registers_reg_19_40_inst : DFF_X1 port map( D => n8471, CK => clk, Q => 
                           n17797, QN => n4063);
   registers_reg_19_39_inst : DFF_X1 port map( D => n8470, CK => clk, Q => 
                           n17796, QN => n4064);
   registers_reg_19_38_inst : DFF_X1 port map( D => n8469, CK => clk, Q => 
                           n17815, QN => n4065);
   registers_reg_19_37_inst : DFF_X1 port map( D => n8468, CK => clk, Q => 
                           n17806, QN => n4066);
   registers_reg_19_36_inst : DFF_X1 port map( D => n8467, CK => clk, Q => 
                           n17805, QN => n4067);
   registers_reg_19_35_inst : DFF_X1 port map( D => n8466, CK => clk, Q => 
                           n17791, QN => n4068);
   registers_reg_19_34_inst : DFF_X1 port map( D => n8465, CK => clk, Q => 
                           n17790, QN => n4069);
   registers_reg_19_33_inst : DFF_X1 port map( D => n8464, CK => clk, Q => 
                           n17789, QN => n4070);
   registers_reg_19_32_inst : DFF_X1 port map( D => n8463, CK => clk, Q => 
                           n17788, QN => n4071);
   registers_reg_19_31_inst : DFF_X1 port map( D => n8462, CK => clk, Q => 
                           n17787, QN => n4072);
   registers_reg_19_30_inst : DFF_X1 port map( D => n8461, CK => clk, Q => 
                           n17786, QN => n4073);
   registers_reg_19_29_inst : DFF_X1 port map( D => n8460, CK => clk, Q => 
                           n17785, QN => n4074);
   registers_reg_19_28_inst : DFF_X1 port map( D => n8459, CK => clk, Q => 
                           n17784, QN => n4075);
   registers_reg_19_27_inst : DFF_X1 port map( D => n8458, CK => clk, Q => 
                           n17783, QN => n4076);
   registers_reg_19_26_inst : DFF_X1 port map( D => n8457, CK => clk, Q => 
                           n17782, QN => n4077);
   registers_reg_19_25_inst : DFF_X1 port map( D => n8456, CK => clk, Q => 
                           n17781, QN => n4078);
   registers_reg_19_24_inst : DFF_X1 port map( D => n8455, CK => clk, Q => 
                           n17780, QN => n4079);
   registers_reg_19_23_inst : DFF_X1 port map( D => n8454, CK => clk, Q => 
                           n17779, QN => n4080);
   registers_reg_19_22_inst : DFF_X1 port map( D => n8453, CK => clk, Q => 
                           n17778, QN => n4081);
   registers_reg_19_21_inst : DFF_X1 port map( D => n8452, CK => clk, Q => 
                           n17777, QN => n4082);
   registers_reg_19_20_inst : DFF_X1 port map( D => n8451, CK => clk, Q => 
                           n17776, QN => n4083);
   registers_reg_19_19_inst : DFF_X1 port map( D => n8450, CK => clk, Q => 
                           n17775, QN => n4084);
   registers_reg_19_18_inst : DFF_X1 port map( D => n8449, CK => clk, Q => 
                           n17774, QN => n4085);
   registers_reg_19_17_inst : DFF_X1 port map( D => n8448, CK => clk, Q => 
                           n17773, QN => n4086);
   registers_reg_19_16_inst : DFF_X1 port map( D => n8447, CK => clk, Q => 
                           n17772, QN => n4087);
   registers_reg_19_15_inst : DFF_X1 port map( D => n8446, CK => clk, Q => 
                           n17771, QN => n4088);
   registers_reg_19_14_inst : DFF_X1 port map( D => n8445, CK => clk, Q => 
                           n17770, QN => n4089);
   registers_reg_19_13_inst : DFF_X1 port map( D => n8444, CK => clk, Q => 
                           n17769, QN => n4090);
   registers_reg_19_12_inst : DFF_X1 port map( D => n8443, CK => clk, Q => 
                           n17768, QN => n4091);
   registers_reg_19_11_inst : DFF_X1 port map( D => n8442, CK => clk, Q => 
                           n17814, QN => n4092);
   registers_reg_19_10_inst : DFF_X1 port map( D => n8441, CK => clk, Q => 
                           n17813, QN => n4093);
   registers_reg_19_9_inst : DFF_X1 port map( D => n8440, CK => clk, Q => 
                           n17812, QN => n4094);
   registers_reg_19_8_inst : DFF_X1 port map( D => n8439, CK => clk, Q => 
                           n17811, QN => n4095);
   registers_reg_19_7_inst : DFF_X1 port map( D => n8438, CK => clk, Q => 
                           n17810, QN => n4096);
   registers_reg_19_6_inst : DFF_X1 port map( D => n8437, CK => clk, Q => 
                           n17809, QN => n4097);
   registers_reg_19_5_inst : DFF_X1 port map( D => n8436, CK => clk, Q => 
                           n17808, QN => n4098);
   registers_reg_19_4_inst : DFF_X1 port map( D => n8435, CK => clk, Q => 
                           n17807, QN => n4099);
   registers_reg_30_54_inst : DFF_X1 port map( D => n9189, CK => clk, Q => 
                           n15859, QN => n3312);
   registers_reg_30_53_inst : DFF_X1 port map( D => n9188, CK => clk, Q => 
                           n15858, QN => n3313);
   registers_reg_30_52_inst : DFF_X1 port map( D => n9187, CK => clk, Q => 
                           n15857, QN => n3314);
   registers_reg_30_51_inst : DFF_X1 port map( D => n9186, CK => clk, Q => 
                           n15856, QN => n3315);
   registers_reg_30_50_inst : DFF_X1 port map( D => n9185, CK => clk, Q => 
                           n15855, QN => n3316);
   registers_reg_30_49_inst : DFF_X1 port map( D => n9184, CK => clk, Q => 
                           n15854, QN => n3317);
   registers_reg_30_48_inst : DFF_X1 port map( D => n9183, CK => clk, Q => 
                           n15853, QN => n3318);
   registers_reg_30_47_inst : DFF_X1 port map( D => n9182, CK => clk, Q => 
                           n15852, QN => n3319);
   registers_reg_30_46_inst : DFF_X1 port map( D => n9181, CK => clk, Q => 
                           n15851, QN => n3320);
   registers_reg_30_45_inst : DFF_X1 port map( D => n9180, CK => clk, Q => 
                           n15850, QN => n3321);
   registers_reg_30_44_inst : DFF_X1 port map( D => n9179, CK => clk, Q => 
                           n15849, QN => n3322);
   registers_reg_30_43_inst : DFF_X1 port map( D => n9178, CK => clk, Q => 
                           n15848, QN => n3323);
   registers_reg_30_42_inst : DFF_X1 port map( D => n9177, CK => clk, Q => 
                           n15847, QN => n3324);
   registers_reg_30_41_inst : DFF_X1 port map( D => n9176, CK => clk, Q => 
                           n15846, QN => n3325);
   registers_reg_30_40_inst : DFF_X1 port map( D => n9175, CK => clk, Q => 
                           n15845, QN => n3326);
   registers_reg_30_39_inst : DFF_X1 port map( D => n9174, CK => clk, Q => 
                           n15844, QN => n3327);
   registers_reg_30_38_inst : DFF_X1 port map( D => n9173, CK => clk, Q => 
                           n15843, QN => n3328);
   registers_reg_30_37_inst : DFF_X1 port map( D => n9172, CK => clk, Q => 
                           n15842, QN => n3329);
   registers_reg_30_36_inst : DFF_X1 port map( D => n9171, CK => clk, Q => 
                           n15841, QN => n3330);
   registers_reg_30_35_inst : DFF_X1 port map( D => n9170, CK => clk, Q => 
                           n15840, QN => n3331);
   registers_reg_30_34_inst : DFF_X1 port map( D => n9169, CK => clk, Q => 
                           n15839, QN => n3332);
   registers_reg_30_33_inst : DFF_X1 port map( D => n9168, CK => clk, Q => 
                           n15838, QN => n3333);
   registers_reg_30_32_inst : DFF_X1 port map( D => n9167, CK => clk, Q => 
                           n15837, QN => n3334);
   registers_reg_30_31_inst : DFF_X1 port map( D => n9166, CK => clk, Q => 
                           n15836, QN => n3335);
   registers_reg_30_30_inst : DFF_X1 port map( D => n9165, CK => clk, Q => 
                           n15835, QN => n3336);
   registers_reg_30_29_inst : DFF_X1 port map( D => n9164, CK => clk, Q => 
                           n15834, QN => n3337);
   registers_reg_30_28_inst : DFF_X1 port map( D => n9163, CK => clk, Q => 
                           n15833, QN => n3338);
   registers_reg_30_27_inst : DFF_X1 port map( D => n9162, CK => clk, Q => 
                           n15832, QN => n3339);
   registers_reg_30_26_inst : DFF_X1 port map( D => n9161, CK => clk, Q => 
                           n15831, QN => n3340);
   registers_reg_30_25_inst : DFF_X1 port map( D => n9160, CK => clk, Q => 
                           n15830, QN => n3341);
   registers_reg_30_24_inst : DFF_X1 port map( D => n9159, CK => clk, Q => 
                           n15829, QN => n3342);
   registers_reg_30_23_inst : DFF_X1 port map( D => n9158, CK => clk, Q => 
                           n15828, QN => n3343);
   registers_reg_30_22_inst : DFF_X1 port map( D => n9157, CK => clk, Q => 
                           n15827, QN => n3344);
   registers_reg_30_21_inst : DFF_X1 port map( D => n9156, CK => clk, Q => 
                           n15826, QN => n3345);
   registers_reg_30_20_inst : DFF_X1 port map( D => n9155, CK => clk, Q => 
                           n15825, QN => n3346);
   registers_reg_30_19_inst : DFF_X1 port map( D => n9154, CK => clk, Q => 
                           n15824, QN => n3347);
   registers_reg_30_18_inst : DFF_X1 port map( D => n9153, CK => clk, Q => 
                           n15823, QN => n3348);
   registers_reg_30_17_inst : DFF_X1 port map( D => n9152, CK => clk, Q => 
                           n15822, QN => n3349);
   registers_reg_30_16_inst : DFF_X1 port map( D => n9151, CK => clk, Q => 
                           n15821, QN => n3350);
   registers_reg_30_15_inst : DFF_X1 port map( D => n9150, CK => clk, Q => 
                           n15820, QN => n3351);
   registers_reg_30_14_inst : DFF_X1 port map( D => n9149, CK => clk, Q => 
                           n15819, QN => n3352);
   registers_reg_30_13_inst : DFF_X1 port map( D => n9148, CK => clk, Q => 
                           n15818, QN => n3353);
   registers_reg_30_12_inst : DFF_X1 port map( D => n9147, CK => clk, Q => 
                           n15817, QN => n3354);
   registers_reg_30_11_inst : DFF_X1 port map( D => n9146, CK => clk, Q => 
                           n15816, QN => n3355);
   registers_reg_30_10_inst : DFF_X1 port map( D => n9145, CK => clk, Q => 
                           n15815, QN => n3356);
   registers_reg_30_9_inst : DFF_X1 port map( D => n9144, CK => clk, Q => 
                           n15814, QN => n3357);
   registers_reg_30_8_inst : DFF_X1 port map( D => n9143, CK => clk, Q => 
                           n15813, QN => n3358);
   registers_reg_30_7_inst : DFF_X1 port map( D => n9142, CK => clk, Q => 
                           n15812, QN => n3359);
   registers_reg_30_6_inst : DFF_X1 port map( D => n9141, CK => clk, Q => 
                           n15811, QN => n3360);
   registers_reg_30_5_inst : DFF_X1 port map( D => n9140, CK => clk, Q => 
                           n15810, QN => n3361);
   registers_reg_30_4_inst : DFF_X1 port map( D => n9139, CK => clk, Q => 
                           n15809, QN => n3362);
   registers_reg_25_63_inst : DFF_X1 port map( D => n8878, CK => clk, Q => 
                           n17700, QN => n3641);
   registers_reg_25_62_inst : DFF_X1 port map( D => n8877, CK => clk, Q => 
                           n17699, QN => n3642);
   registers_reg_25_61_inst : DFF_X1 port map( D => n8876, CK => clk, Q => 
                           n17698, QN => n3643);
   registers_reg_25_60_inst : DFF_X1 port map( D => n8875, CK => clk, Q => 
                           n17697, QN => n3644);
   registers_reg_25_59_inst : DFF_X1 port map( D => n8874, CK => clk, Q => 
                           n17721, QN => n3645);
   registers_reg_25_58_inst : DFF_X1 port map( D => n8873, CK => clk, Q => 
                           n17720, QN => n3646);
   registers_reg_25_57_inst : DFF_X1 port map( D => n8872, CK => clk, Q => 
                           n17719, QN => n3647);
   registers_reg_25_56_inst : DFF_X1 port map( D => n8871, CK => clk, Q => 
                           n17718, QN => n3648);
   registers_reg_25_55_inst : DFF_X1 port map( D => n8870, CK => clk, Q => 
                           n17717, QN => n3649);
   registers_reg_25_54_inst : DFF_X1 port map( D => n8869, CK => clk, Q => 
                           n17716, QN => n3650);
   registers_reg_25_53_inst : DFF_X1 port map( D => n8868, CK => clk, Q => 
                           n17715, QN => n3651);
   registers_reg_25_52_inst : DFF_X1 port map( D => n8867, CK => clk, Q => 
                           n17714, QN => n3652);
   registers_reg_25_51_inst : DFF_X1 port map( D => n8866, CK => clk, Q => 
                           n17713, QN => n3653);
   registers_reg_25_50_inst : DFF_X1 port map( D => n8865, CK => clk, Q => 
                           n17712, QN => n3654);
   registers_reg_25_49_inst : DFF_X1 port map( D => n8864, CK => clk, Q => 
                           n17711, QN => n3655);
   registers_reg_25_48_inst : DFF_X1 port map( D => n8863, CK => clk, Q => 
                           n17710, QN => n3656);
   registers_reg_25_47_inst : DFF_X1 port map( D => n8862, CK => clk, Q => 
                           n17709, QN => n3657);
   registers_reg_25_46_inst : DFF_X1 port map( D => n8861, CK => clk, Q => 
                           n17708, QN => n3658);
   registers_reg_25_45_inst : DFF_X1 port map( D => n8860, CK => clk, Q => 
                           n17707, QN => n3659);
   registers_reg_25_44_inst : DFF_X1 port map( D => n8859, CK => clk, Q => 
                           n17706, QN => n3660);
   registers_reg_25_43_inst : DFF_X1 port map( D => n8858, CK => clk, Q => 
                           n17705, QN => n3661);
   registers_reg_25_42_inst : DFF_X1 port map( D => n8857, CK => clk, Q => 
                           n17704, QN => n3662);
   registers_reg_25_41_inst : DFF_X1 port map( D => n8856, CK => clk, Q => 
                           n17703, QN => n3663);
   registers_reg_25_40_inst : DFF_X1 port map( D => n8855, CK => clk, Q => 
                           n17702, QN => n3664);
   registers_reg_25_39_inst : DFF_X1 port map( D => n8854, CK => clk, Q => 
                           n17701, QN => n3665);
   registers_reg_25_38_inst : DFF_X1 port map( D => n8853, CK => clk, Q => 
                           n17696, QN => n3666);
   registers_reg_25_37_inst : DFF_X1 port map( D => n8852, CK => clk, Q => 
                           n17755, QN => n3667);
   registers_reg_25_36_inst : DFF_X1 port map( D => n8851, CK => clk, Q => 
                           n17754, QN => n3668);
   registers_reg_25_35_inst : DFF_X1 port map( D => n8850, CK => clk, Q => 
                           n17753, QN => n3669);
   registers_reg_25_34_inst : DFF_X1 port map( D => n8849, CK => clk, Q => 
                           n17752, QN => n3670);
   registers_reg_25_33_inst : DFF_X1 port map( D => n8848, CK => clk, Q => 
                           n17751, QN => n3671);
   registers_reg_25_32_inst : DFF_X1 port map( D => n8847, CK => clk, Q => 
                           n17750, QN => n3672);
   registers_reg_25_31_inst : DFF_X1 port map( D => n8846, CK => clk, Q => 
                           n17749, QN => n3673);
   registers_reg_25_30_inst : DFF_X1 port map( D => n8845, CK => clk, Q => 
                           n17748, QN => n3674);
   registers_reg_25_29_inst : DFF_X1 port map( D => n8844, CK => clk, Q => 
                           n17747, QN => n3675);
   registers_reg_25_28_inst : DFF_X1 port map( D => n8843, CK => clk, Q => 
                           n17746, QN => n3676);
   registers_reg_25_27_inst : DFF_X1 port map( D => n8842, CK => clk, Q => 
                           n17745, QN => n3677);
   registers_reg_25_26_inst : DFF_X1 port map( D => n8841, CK => clk, Q => 
                           n17744, QN => n3678);
   registers_reg_25_25_inst : DFF_X1 port map( D => n8840, CK => clk, Q => 
                           n17743, QN => n3679);
   registers_reg_25_24_inst : DFF_X1 port map( D => n8839, CK => clk, Q => 
                           n17742, QN => n3680);
   registers_reg_25_23_inst : DFF_X1 port map( D => n8838, CK => clk, Q => 
                           n17741, QN => n3681);
   registers_reg_25_22_inst : DFF_X1 port map( D => n8837, CK => clk, Q => 
                           n17740, QN => n3682);
   registers_reg_25_21_inst : DFF_X1 port map( D => n8836, CK => clk, Q => 
                           n17739, QN => n3683);
   registers_reg_25_20_inst : DFF_X1 port map( D => n8835, CK => clk, Q => 
                           n17738, QN => n3684);
   registers_reg_25_19_inst : DFF_X1 port map( D => n8834, CK => clk, Q => 
                           n17737, QN => n3685);
   registers_reg_25_18_inst : DFF_X1 port map( D => n8833, CK => clk, Q => 
                           n17736, QN => n3686);
   registers_reg_25_17_inst : DFF_X1 port map( D => n8832, CK => clk, Q => 
                           n17735, QN => n3687);
   registers_reg_25_16_inst : DFF_X1 port map( D => n8831, CK => clk, Q => 
                           n17734, QN => n3688);
   registers_reg_25_15_inst : DFF_X1 port map( D => n8830, CK => clk, Q => 
                           n17733, QN => n3689);
   registers_reg_25_14_inst : DFF_X1 port map( D => n8829, CK => clk, Q => 
                           n17732, QN => n3690);
   registers_reg_25_13_inst : DFF_X1 port map( D => n8828, CK => clk, Q => 
                           n17731, QN => n3691);
   registers_reg_25_12_inst : DFF_X1 port map( D => n8827, CK => clk, Q => 
                           n17730, QN => n3692);
   registers_reg_25_11_inst : DFF_X1 port map( D => n8826, CK => clk, Q => 
                           n17729, QN => n3693);
   registers_reg_25_10_inst : DFF_X1 port map( D => n8825, CK => clk, Q => 
                           n17728, QN => n3694);
   registers_reg_25_9_inst : DFF_X1 port map( D => n8824, CK => clk, Q => 
                           n17727, QN => n3695);
   registers_reg_25_8_inst : DFF_X1 port map( D => n8823, CK => clk, Q => 
                           n17726, QN => n3696);
   registers_reg_25_7_inst : DFF_X1 port map( D => n8822, CK => clk, Q => 
                           n17725, QN => n3697);
   registers_reg_25_6_inst : DFF_X1 port map( D => n8821, CK => clk, Q => 
                           n17724, QN => n3698);
   registers_reg_25_5_inst : DFF_X1 port map( D => n8820, CK => clk, Q => 
                           n17723, QN => n3699);
   registers_reg_25_4_inst : DFF_X1 port map( D => n8819, CK => clk, Q => 
                           n17722, QN => n3700);
   registers_reg_24_63_inst : DFF_X1 port map( D => n8814, CK => clk, Q => 
                           n17867, QN => n3707);
   registers_reg_24_62_inst : DFF_X1 port map( D => n8813, CK => clk, Q => 
                           n17866, QN => n3708);
   registers_reg_24_61_inst : DFF_X1 port map( D => n8812, CK => clk, Q => 
                           n17865, QN => n3709);
   registers_reg_24_60_inst : DFF_X1 port map( D => n8811, CK => clk, Q => 
                           n17864, QN => n3710);
   registers_reg_24_59_inst : DFF_X1 port map( D => n8810, CK => clk, Q => 
                           n17863, QN => n3711);
   registers_reg_24_58_inst : DFF_X1 port map( D => n8809, CK => clk, Q => 
                           n17862, QN => n3712);
   registers_reg_24_57_inst : DFF_X1 port map( D => n8808, CK => clk, Q => 
                           n17861, QN => n3713);
   registers_reg_24_56_inst : DFF_X1 port map( D => n8807, CK => clk, Q => 
                           n17860, QN => n3714);
   registers_reg_24_55_inst : DFF_X1 port map( D => n8806, CK => clk, Q => 
                           n17859, QN => n3715);
   registers_reg_24_54_inst : DFF_X1 port map( D => n8805, CK => clk, Q => 
                           n17858, QN => n3716);
   registers_reg_24_53_inst : DFF_X1 port map( D => n8804, CK => clk, Q => 
                           n17857, QN => n3717);
   registers_reg_24_52_inst : DFF_X1 port map( D => n8803, CK => clk, Q => 
                           n17856, QN => n3718);
   registers_reg_24_51_inst : DFF_X1 port map( D => n8802, CK => clk, Q => 
                           n17855, QN => n3719);
   registers_reg_24_50_inst : DFF_X1 port map( D => n8801, CK => clk, Q => 
                           n17854, QN => n3720);
   registers_reg_24_49_inst : DFF_X1 port map( D => n8800, CK => clk, Q => 
                           n17853, QN => n3721);
   registers_reg_24_48_inst : DFF_X1 port map( D => n8799, CK => clk, Q => 
                           n17852, QN => n3722);
   registers_reg_24_47_inst : DFF_X1 port map( D => n8798, CK => clk, Q => 
                           n17851, QN => n3723);
   registers_reg_24_46_inst : DFF_X1 port map( D => n8797, CK => clk, Q => 
                           n17850, QN => n3724);
   registers_reg_24_45_inst : DFF_X1 port map( D => n8796, CK => clk, Q => 
                           n17849, QN => n3725);
   registers_reg_24_44_inst : DFF_X1 port map( D => n8795, CK => clk, Q => 
                           n17848, QN => n3726);
   registers_reg_24_43_inst : DFF_X1 port map( D => n8794, CK => clk, Q => 
                           n17847, QN => n3727);
   registers_reg_24_42_inst : DFF_X1 port map( D => n8793, CK => clk, Q => 
                           n17846, QN => n3728);
   registers_reg_24_41_inst : DFF_X1 port map( D => n8792, CK => clk, Q => 
                           n17845, QN => n3729);
   registers_reg_24_40_inst : DFF_X1 port map( D => n8791, CK => clk, Q => 
                           n17844, QN => n3730);
   registers_reg_24_39_inst : DFF_X1 port map( D => n8790, CK => clk, Q => 
                           n17843, QN => n3731);
   registers_reg_24_38_inst : DFF_X1 port map( D => n8789, CK => clk, Q => 
                           n17842, QN => n3732);
   registers_reg_24_37_inst : DFF_X1 port map( D => n8788, CK => clk, Q => 
                           n17841, QN => n3733);
   registers_reg_24_36_inst : DFF_X1 port map( D => n8787, CK => clk, Q => 
                           n17840, QN => n3734);
   registers_reg_24_35_inst : DFF_X1 port map( D => n8786, CK => clk, Q => 
                           n17839, QN => n3735);
   registers_reg_24_34_inst : DFF_X1 port map( D => n8785, CK => clk, Q => 
                           n17838, QN => n3736);
   registers_reg_24_33_inst : DFF_X1 port map( D => n8784, CK => clk, Q => 
                           n17837, QN => n3737);
   registers_reg_24_32_inst : DFF_X1 port map( D => n8783, CK => clk, Q => 
                           n17836, QN => n3738);
   registers_reg_24_31_inst : DFF_X1 port map( D => n8782, CK => clk, Q => 
                           n17835, QN => n3739);
   registers_reg_24_30_inst : DFF_X1 port map( D => n8781, CK => clk, Q => 
                           n17834, QN => n3740);
   registers_reg_24_29_inst : DFF_X1 port map( D => n8780, CK => clk, Q => 
                           n17833, QN => n3741);
   registers_reg_24_28_inst : DFF_X1 port map( D => n8779, CK => clk, Q => 
                           n17832, QN => n3742);
   registers_reg_24_27_inst : DFF_X1 port map( D => n8778, CK => clk, Q => 
                           n17831, QN => n3743);
   registers_reg_24_26_inst : DFF_X1 port map( D => n8777, CK => clk, Q => 
                           n17830, QN => n3744);
   registers_reg_24_25_inst : DFF_X1 port map( D => n8776, CK => clk, Q => 
                           n17829, QN => n3745);
   registers_reg_24_24_inst : DFF_X1 port map( D => n8775, CK => clk, Q => 
                           n17828, QN => n3746);
   registers_reg_24_23_inst : DFF_X1 port map( D => n8774, CK => clk, Q => 
                           n17827, QN => n3747);
   registers_reg_24_22_inst : DFF_X1 port map( D => n8773, CK => clk, Q => 
                           n17826, QN => n3748);
   registers_reg_24_21_inst : DFF_X1 port map( D => n8772, CK => clk, Q => 
                           n17825, QN => n3749);
   registers_reg_24_20_inst : DFF_X1 port map( D => n8771, CK => clk, Q => 
                           n17824, QN => n3750);
   registers_reg_24_19_inst : DFF_X1 port map( D => n8770, CK => clk, Q => 
                           n17823, QN => n3751);
   registers_reg_24_18_inst : DFF_X1 port map( D => n8769, CK => clk, Q => 
                           n17822, QN => n3752);
   registers_reg_24_17_inst : DFF_X1 port map( D => n8768, CK => clk, Q => 
                           n17821, QN => n3753);
   registers_reg_24_16_inst : DFF_X1 port map( D => n8767, CK => clk, Q => 
                           n17820, QN => n3754);
   registers_reg_24_15_inst : DFF_X1 port map( D => n8766, CK => clk, Q => 
                           n17819, QN => n3755);
   registers_reg_24_14_inst : DFF_X1 port map( D => n8765, CK => clk, Q => 
                           n17818, QN => n3756);
   registers_reg_24_13_inst : DFF_X1 port map( D => n8764, CK => clk, Q => 
                           n17817, QN => n3757);
   registers_reg_24_12_inst : DFF_X1 port map( D => n8763, CK => clk, Q => 
                           n17816, QN => n3758);
   registers_reg_24_11_inst : DFF_X1 port map( D => n8762, CK => clk, Q => 
                           n17875, QN => n3759);
   registers_reg_24_10_inst : DFF_X1 port map( D => n8761, CK => clk, Q => 
                           n17874, QN => n3760);
   registers_reg_24_9_inst : DFF_X1 port map( D => n8760, CK => clk, Q => 
                           n17873, QN => n3761);
   registers_reg_24_8_inst : DFF_X1 port map( D => n8759, CK => clk, Q => 
                           n17872, QN => n3762);
   registers_reg_24_7_inst : DFF_X1 port map( D => n8758, CK => clk, Q => 
                           n17871, QN => n3763);
   registers_reg_24_6_inst : DFF_X1 port map( D => n8757, CK => clk, Q => 
                           n17870, QN => n3764);
   registers_reg_24_5_inst : DFF_X1 port map( D => n8756, CK => clk, Q => 
                           n17869, QN => n3765);
   registers_reg_24_4_inst : DFF_X1 port map( D => n8755, CK => clk, Q => 
                           n17868, QN => n3766);
   registers_reg_17_63_inst : DFF_X1 port map( D => n8366, CK => clk, Q => 
                           n15476, QN => n4179);
   registers_reg_17_62_inst : DFF_X1 port map( D => n8365, CK => clk, Q => 
                           n15475, QN => n4180);
   registers_reg_17_61_inst : DFF_X1 port map( D => n8364, CK => clk, Q => 
                           n15474, QN => n4181);
   registers_reg_17_60_inst : DFF_X1 port map( D => n8363, CK => clk, Q => 
                           n15473, QN => n4182);
   registers_reg_17_59_inst : DFF_X1 port map( D => n8362, CK => clk, Q => 
                           n15472, QN => n4183);
   registers_reg_17_58_inst : DFF_X1 port map( D => n8361, CK => clk, Q => 
                           n15471, QN => n4184);
   registers_reg_17_57_inst : DFF_X1 port map( D => n8360, CK => clk, Q => 
                           n15470, QN => n4185);
   registers_reg_17_56_inst : DFF_X1 port map( D => n8359, CK => clk, Q => 
                           n15469, QN => n4186);
   registers_reg_17_55_inst : DFF_X1 port map( D => n8358, CK => clk, Q => 
                           n15468, QN => n4187);
   registers_reg_17_54_inst : DFF_X1 port map( D => n8357, CK => clk, Q => 
                           n15467, QN => n4188);
   registers_reg_17_53_inst : DFF_X1 port map( D => n8356, CK => clk, Q => 
                           n15466, QN => n4189);
   registers_reg_17_52_inst : DFF_X1 port map( D => n8355, CK => clk, Q => 
                           n15465, QN => n4190);
   registers_reg_17_51_inst : DFF_X1 port map( D => n8354, CK => clk, Q => 
                           n15464, QN => n4191);
   registers_reg_17_50_inst : DFF_X1 port map( D => n8353, CK => clk, Q => 
                           n15463, QN => n4192);
   registers_reg_17_49_inst : DFF_X1 port map( D => n8352, CK => clk, Q => 
                           n15462, QN => n4193);
   registers_reg_17_48_inst : DFF_X1 port map( D => n8351, CK => clk, Q => 
                           n15461, QN => n4194);
   registers_reg_17_47_inst : DFF_X1 port map( D => n8350, CK => clk, Q => 
                           n15460, QN => n4195);
   registers_reg_17_46_inst : DFF_X1 port map( D => n8349, CK => clk, Q => 
                           n15459, QN => n4196);
   registers_reg_17_45_inst : DFF_X1 port map( D => n8348, CK => clk, Q => 
                           n15458, QN => n4197);
   registers_reg_17_44_inst : DFF_X1 port map( D => n8347, CK => clk, Q => 
                           n15457, QN => n4198);
   registers_reg_17_43_inst : DFF_X1 port map( D => n8346, CK => clk, Q => 
                           n15456, QN => n4199);
   registers_reg_17_42_inst : DFF_X1 port map( D => n8345, CK => clk, Q => 
                           n15455, QN => n4200);
   registers_reg_17_41_inst : DFF_X1 port map( D => n8344, CK => clk, Q => 
                           n15454, QN => n4201);
   registers_reg_17_40_inst : DFF_X1 port map( D => n8343, CK => clk, Q => 
                           n15453, QN => n4202);
   registers_reg_17_39_inst : DFF_X1 port map( D => n8342, CK => clk, Q => 
                           n15452, QN => n4203);
   registers_reg_17_38_inst : DFF_X1 port map( D => n8341, CK => clk, Q => 
                           n15451, QN => n4204);
   registers_reg_17_37_inst : DFF_X1 port map( D => n8340, CK => clk, Q => 
                           n15450, QN => n4205);
   registers_reg_17_36_inst : DFF_X1 port map( D => n8339, CK => clk, Q => 
                           n15449, QN => n4206);
   registers_reg_17_35_inst : DFF_X1 port map( D => n8338, CK => clk, Q => 
                           n15448, QN => n4207);
   registers_reg_17_34_inst : DFF_X1 port map( D => n8337, CK => clk, Q => 
                           n15447, QN => n4208);
   registers_reg_17_33_inst : DFF_X1 port map( D => n8336, CK => clk, Q => 
                           n15446, QN => n4209);
   registers_reg_17_32_inst : DFF_X1 port map( D => n8335, CK => clk, Q => 
                           n15445, QN => n4210);
   registers_reg_17_31_inst : DFF_X1 port map( D => n8334, CK => clk, Q => 
                           n15444, QN => n4211);
   registers_reg_17_30_inst : DFF_X1 port map( D => n8333, CK => clk, Q => 
                           n15443, QN => n4212);
   registers_reg_17_29_inst : DFF_X1 port map( D => n8332, CK => clk, Q => 
                           n15442, QN => n4213);
   registers_reg_17_28_inst : DFF_X1 port map( D => n8331, CK => clk, Q => 
                           n15441, QN => n4214);
   registers_reg_17_27_inst : DFF_X1 port map( D => n8330, CK => clk, Q => 
                           n15440, QN => n4215);
   registers_reg_17_26_inst : DFF_X1 port map( D => n8329, CK => clk, Q => 
                           n15439, QN => n4216);
   registers_reg_17_25_inst : DFF_X1 port map( D => n8328, CK => clk, Q => 
                           n15438, QN => n4217);
   registers_reg_17_24_inst : DFF_X1 port map( D => n8327, CK => clk, Q => 
                           n15437, QN => n4218);
   registers_reg_17_23_inst : DFF_X1 port map( D => n8326, CK => clk, Q => 
                           n15436, QN => n4219);
   registers_reg_17_22_inst : DFF_X1 port map( D => n8325, CK => clk, Q => 
                           n15435, QN => n4220);
   registers_reg_17_21_inst : DFF_X1 port map( D => n8324, CK => clk, Q => 
                           n15434, QN => n4221);
   registers_reg_17_20_inst : DFF_X1 port map( D => n8323, CK => clk, Q => 
                           n15433, QN => n4222);
   registers_reg_17_19_inst : DFF_X1 port map( D => n8322, CK => clk, Q => 
                           n15432, QN => n4223);
   registers_reg_17_18_inst : DFF_X1 port map( D => n8321, CK => clk, Q => 
                           n15431, QN => n4224);
   registers_reg_17_17_inst : DFF_X1 port map( D => n8320, CK => clk, Q => 
                           n15430, QN => n4225);
   registers_reg_17_16_inst : DFF_X1 port map( D => n8319, CK => clk, Q => 
                           n15429, QN => n4226);
   registers_reg_17_15_inst : DFF_X1 port map( D => n8318, CK => clk, Q => 
                           n15428, QN => n4227);
   registers_reg_17_14_inst : DFF_X1 port map( D => n8317, CK => clk, Q => 
                           n15427, QN => n4228);
   registers_reg_17_13_inst : DFF_X1 port map( D => n8316, CK => clk, Q => 
                           n15426, QN => n4229);
   registers_reg_17_12_inst : DFF_X1 port map( D => n8315, CK => clk, Q => 
                           n15425, QN => n4230);
   registers_reg_17_11_inst : DFF_X1 port map( D => n8314, CK => clk, Q => 
                           n15424, QN => n4231);
   registers_reg_17_10_inst : DFF_X1 port map( D => n8313, CK => clk, Q => 
                           n15423, QN => n4232);
   registers_reg_17_9_inst : DFF_X1 port map( D => n8312, CK => clk, Q => 
                           n15422, QN => n4233);
   registers_reg_17_8_inst : DFF_X1 port map( D => n8311, CK => clk, Q => 
                           n15421, QN => n4234);
   registers_reg_17_7_inst : DFF_X1 port map( D => n8310, CK => clk, Q => 
                           n15420, QN => n4235);
   registers_reg_17_6_inst : DFF_X1 port map( D => n8309, CK => clk, Q => 
                           n15419, QN => n4236);
   registers_reg_17_5_inst : DFF_X1 port map( D => n8308, CK => clk, Q => 
                           n15418, QN => n4237);
   registers_reg_17_4_inst : DFF_X1 port map( D => n8307, CK => clk, Q => 
                           n15417, QN => n4238);
   registers_reg_29_63_inst : DFF_X1 port map( D => n9134, CK => clk, Q => 
                           n15356, QN => n3371);
   registers_reg_29_62_inst : DFF_X1 port map( D => n9133, CK => clk, Q => 
                           n15355, QN => n3372);
   registers_reg_29_61_inst : DFF_X1 port map( D => n9132, CK => clk, Q => 
                           n15354, QN => n3373);
   registers_reg_29_60_inst : DFF_X1 port map( D => n9131, CK => clk, Q => 
                           n15353, QN => n3374);
   registers_reg_29_59_inst : DFF_X1 port map( D => n9130, CK => clk, Q => 
                           n15352, QN => n3375);
   registers_reg_29_58_inst : DFF_X1 port map( D => n9129, CK => clk, Q => 
                           n15351, QN => n3376);
   registers_reg_29_57_inst : DFF_X1 port map( D => n9128, CK => clk, Q => 
                           n15350, QN => n3377);
   registers_reg_29_56_inst : DFF_X1 port map( D => n9127, CK => clk, Q => 
                           n15349, QN => n3378);
   registers_reg_29_55_inst : DFF_X1 port map( D => n9126, CK => clk, Q => 
                           n15348, QN => n3379);
   registers_reg_29_54_inst : DFF_X1 port map( D => n9125, CK => clk, Q => 
                           n15347, QN => n3380);
   registers_reg_29_53_inst : DFF_X1 port map( D => n9124, CK => clk, Q => 
                           n15346, QN => n3381);
   registers_reg_29_52_inst : DFF_X1 port map( D => n9123, CK => clk, Q => 
                           n15345, QN => n3382);
   registers_reg_29_51_inst : DFF_X1 port map( D => n9122, CK => clk, Q => 
                           n15344, QN => n3383);
   registers_reg_29_50_inst : DFF_X1 port map( D => n9121, CK => clk, Q => 
                           n15343, QN => n3384);
   registers_reg_29_49_inst : DFF_X1 port map( D => n9120, CK => clk, Q => 
                           n15342, QN => n3385);
   registers_reg_29_48_inst : DFF_X1 port map( D => n9119, CK => clk, Q => 
                           n15341, QN => n3386);
   registers_reg_29_47_inst : DFF_X1 port map( D => n9118, CK => clk, Q => 
                           n15340, QN => n3387);
   registers_reg_29_46_inst : DFF_X1 port map( D => n9117, CK => clk, Q => 
                           n15339, QN => n3388);
   registers_reg_29_45_inst : DFF_X1 port map( D => n9116, CK => clk, Q => 
                           n15338, QN => n3389);
   registers_reg_29_44_inst : DFF_X1 port map( D => n9115, CK => clk, Q => 
                           n15337, QN => n3390);
   registers_reg_29_43_inst : DFF_X1 port map( D => n9114, CK => clk, Q => 
                           n15336, QN => n3391);
   registers_reg_29_42_inst : DFF_X1 port map( D => n9113, CK => clk, Q => 
                           n15335, QN => n3392);
   registers_reg_29_41_inst : DFF_X1 port map( D => n9112, CK => clk, Q => 
                           n15334, QN => n3393);
   registers_reg_29_40_inst : DFF_X1 port map( D => n9111, CK => clk, Q => 
                           n15333, QN => n3394);
   registers_reg_29_39_inst : DFF_X1 port map( D => n9110, CK => clk, Q => 
                           n15332, QN => n3395);
   registers_reg_29_38_inst : DFF_X1 port map( D => n9109, CK => clk, Q => 
                           n15331, QN => n3396);
   registers_reg_29_37_inst : DFF_X1 port map( D => n9108, CK => clk, Q => 
                           n15330, QN => n3397);
   registers_reg_29_36_inst : DFF_X1 port map( D => n9107, CK => clk, Q => 
                           n15329, QN => n3398);
   registers_reg_29_35_inst : DFF_X1 port map( D => n9106, CK => clk, Q => 
                           n15328, QN => n3399);
   registers_reg_29_34_inst : DFF_X1 port map( D => n9105, CK => clk, Q => 
                           n15327, QN => n3400);
   registers_reg_29_33_inst : DFF_X1 port map( D => n9104, CK => clk, Q => 
                           n15326, QN => n3401);
   registers_reg_29_32_inst : DFF_X1 port map( D => n9103, CK => clk, Q => 
                           n15325, QN => n3402);
   registers_reg_29_31_inst : DFF_X1 port map( D => n9102, CK => clk, Q => 
                           n15324, QN => n3403);
   registers_reg_29_30_inst : DFF_X1 port map( D => n9101, CK => clk, Q => 
                           n15323, QN => n3404);
   registers_reg_29_29_inst : DFF_X1 port map( D => n9100, CK => clk, Q => 
                           n15322, QN => n3405);
   registers_reg_29_28_inst : DFF_X1 port map( D => n9099, CK => clk, Q => 
                           n15321, QN => n3406);
   registers_reg_29_27_inst : DFF_X1 port map( D => n9098, CK => clk, Q => 
                           n15320, QN => n3407);
   registers_reg_29_26_inst : DFF_X1 port map( D => n9097, CK => clk, Q => 
                           n15319, QN => n3408);
   registers_reg_29_25_inst : DFF_X1 port map( D => n9096, CK => clk, Q => 
                           n15318, QN => n3409);
   registers_reg_29_24_inst : DFF_X1 port map( D => n9095, CK => clk, Q => 
                           n15317, QN => n3410);
   registers_reg_29_23_inst : DFF_X1 port map( D => n9094, CK => clk, Q => 
                           n15316, QN => n3411);
   registers_reg_29_22_inst : DFF_X1 port map( D => n9093, CK => clk, Q => 
                           n15315, QN => n3412);
   registers_reg_29_21_inst : DFF_X1 port map( D => n9092, CK => clk, Q => 
                           n15314, QN => n3413);
   registers_reg_29_20_inst : DFF_X1 port map( D => n9091, CK => clk, Q => 
                           n15313, QN => n3414);
   registers_reg_29_19_inst : DFF_X1 port map( D => n9090, CK => clk, Q => 
                           n15312, QN => n3415);
   registers_reg_29_18_inst : DFF_X1 port map( D => n9089, CK => clk, Q => 
                           n15311, QN => n3416);
   registers_reg_29_17_inst : DFF_X1 port map( D => n9088, CK => clk, Q => 
                           n15310, QN => n3417);
   registers_reg_29_16_inst : DFF_X1 port map( D => n9087, CK => clk, Q => 
                           n15309, QN => n3418);
   registers_reg_29_15_inst : DFF_X1 port map( D => n9086, CK => clk, Q => 
                           n15308, QN => n3419);
   registers_reg_29_14_inst : DFF_X1 port map( D => n9085, CK => clk, Q => 
                           n15307, QN => n3420);
   registers_reg_29_13_inst : DFF_X1 port map( D => n9084, CK => clk, Q => 
                           n15306, QN => n3421);
   registers_reg_29_12_inst : DFF_X1 port map( D => n9083, CK => clk, Q => 
                           n15305, QN => n3422);
   registers_reg_29_11_inst : DFF_X1 port map( D => n9082, CK => clk, Q => 
                           n15304, QN => n3423);
   registers_reg_29_10_inst : DFF_X1 port map( D => n9081, CK => clk, Q => 
                           n15303, QN => n3424);
   registers_reg_29_9_inst : DFF_X1 port map( D => n9080, CK => clk, Q => 
                           n15302, QN => n3425);
   registers_reg_29_8_inst : DFF_X1 port map( D => n9079, CK => clk, Q => 
                           n15301, QN => n3426);
   registers_reg_29_7_inst : DFF_X1 port map( D => n9078, CK => clk, Q => 
                           n15300, QN => n3427);
   registers_reg_29_6_inst : DFF_X1 port map( D => n9077, CK => clk, Q => 
                           n15299, QN => n3428);
   registers_reg_29_5_inst : DFF_X1 port map( D => n9076, CK => clk, Q => 
                           n15298, QN => n3429);
   registers_reg_29_4_inst : DFF_X1 port map( D => n9075, CK => clk, Q => 
                           n15297, QN => n3430);
   registers_reg_5_63_inst : DFF_X1 port map( D => n7598, CK => clk, Q => 
                           n17995, QN => n4990);
   registers_reg_5_62_inst : DFF_X1 port map( D => n7597, CK => clk, Q => 
                           n17994, QN => n4991);
   registers_reg_5_61_inst : DFF_X1 port map( D => n7596, CK => clk, Q => 
                           n17993, QN => n4992);
   registers_reg_5_60_inst : DFF_X1 port map( D => n7595, CK => clk, Q => 
                           n17992, QN => n4993);
   registers_reg_5_59_inst : DFF_X1 port map( D => n7594, CK => clk, Q => 
                           n17991, QN => n4994);
   registers_reg_5_58_inst : DFF_X1 port map( D => n7593, CK => clk, Q => 
                           n17990, QN => n4995);
   registers_reg_5_57_inst : DFF_X1 port map( D => n7592, CK => clk, Q => 
                           n17989, QN => n4996);
   registers_reg_5_56_inst : DFF_X1 port map( D => n7591, CK => clk, Q => 
                           n17988, QN => n4997);
   registers_reg_5_55_inst : DFF_X1 port map( D => n7590, CK => clk, Q => 
                           n17987, QN => n4998);
   registers_reg_5_54_inst : DFF_X1 port map( D => n7589, CK => clk, Q => 
                           n17986, QN => n4999);
   registers_reg_5_53_inst : DFF_X1 port map( D => n7588, CK => clk, Q => 
                           n17985, QN => n5000);
   registers_reg_5_52_inst : DFF_X1 port map( D => n7587, CK => clk, Q => 
                           n17984, QN => n5001);
   registers_reg_5_51_inst : DFF_X1 port map( D => n7586, CK => clk, Q => 
                           n17983, QN => n5002);
   registers_reg_5_50_inst : DFF_X1 port map( D => n7585, CK => clk, Q => 
                           n17982, QN => n5003);
   registers_reg_5_49_inst : DFF_X1 port map( D => n7584, CK => clk, Q => 
                           n17981, QN => n5004);
   registers_reg_5_48_inst : DFF_X1 port map( D => n7583, CK => clk, Q => 
                           n17980, QN => n5005);
   registers_reg_5_47_inst : DFF_X1 port map( D => n7582, CK => clk, Q => 
                           n17979, QN => n5006);
   registers_reg_5_46_inst : DFF_X1 port map( D => n7581, CK => clk, Q => 
                           n17978, QN => n5007);
   registers_reg_5_45_inst : DFF_X1 port map( D => n7580, CK => clk, Q => 
                           n17977, QN => n5008);
   registers_reg_5_44_inst : DFF_X1 port map( D => n7579, CK => clk, Q => 
                           n17976, QN => n5009);
   registers_reg_5_43_inst : DFF_X1 port map( D => n7578, CK => clk, Q => 
                           n17975, QN => n5010);
   registers_reg_5_42_inst : DFF_X1 port map( D => n7577, CK => clk, Q => 
                           n17974, QN => n5011);
   registers_reg_5_41_inst : DFF_X1 port map( D => n7576, CK => clk, Q => 
                           n17973, QN => n5012);
   registers_reg_5_40_inst : DFF_X1 port map( D => n7575, CK => clk, Q => 
                           n17972, QN => n5013);
   registers_reg_5_39_inst : DFF_X1 port map( D => n7574, CK => clk, Q => 
                           n17971, QN => n5014);
   registers_reg_5_38_inst : DFF_X1 port map( D => n7573, CK => clk, Q => 
                           n17970, QN => n5015);
   registers_reg_5_37_inst : DFF_X1 port map( D => n7572, CK => clk, Q => 
                           n17969, QN => n5016);
   registers_reg_5_36_inst : DFF_X1 port map( D => n7571, CK => clk, Q => 
                           n17968, QN => n5017);
   registers_reg_5_35_inst : DFF_X1 port map( D => n7570, CK => clk, Q => 
                           n17967, QN => n5018);
   registers_reg_5_34_inst : DFF_X1 port map( D => n7569, CK => clk, Q => 
                           n17966, QN => n5019);
   registers_reg_5_33_inst : DFF_X1 port map( D => n7568, CK => clk, Q => 
                           n17965, QN => n5020);
   registers_reg_5_32_inst : DFF_X1 port map( D => n7567, CK => clk, Q => 
                           n17964, QN => n5021);
   registers_reg_5_31_inst : DFF_X1 port map( D => n7566, CK => clk, Q => 
                           n17963, QN => n5022);
   registers_reg_5_30_inst : DFF_X1 port map( D => n7565, CK => clk, Q => 
                           n17962, QN => n5023);
   registers_reg_5_29_inst : DFF_X1 port map( D => n7564, CK => clk, Q => 
                           n17961, QN => n5024);
   registers_reg_5_28_inst : DFF_X1 port map( D => n7563, CK => clk, Q => 
                           n17960, QN => n5025);
   registers_reg_5_27_inst : DFF_X1 port map( D => n7562, CK => clk, Q => 
                           n17959, QN => n5026);
   registers_reg_5_26_inst : DFF_X1 port map( D => n7561, CK => clk, Q => 
                           n17958, QN => n5027);
   registers_reg_5_25_inst : DFF_X1 port map( D => n7560, CK => clk, Q => 
                           n17957, QN => n5028);
   registers_reg_5_24_inst : DFF_X1 port map( D => n7559, CK => clk, Q => 
                           n17956, QN => n5029);
   registers_reg_5_23_inst : DFF_X1 port map( D => n7558, CK => clk, Q => 
                           n17955, QN => n5030);
   registers_reg_5_22_inst : DFF_X1 port map( D => n7557, CK => clk, Q => 
                           n17954, QN => n5031);
   registers_reg_5_21_inst : DFF_X1 port map( D => n7556, CK => clk, Q => 
                           n17953, QN => n5032);
   registers_reg_5_20_inst : DFF_X1 port map( D => n7555, CK => clk, Q => 
                           n17952, QN => n5033);
   registers_reg_5_19_inst : DFF_X1 port map( D => n7554, CK => clk, Q => 
                           n17951, QN => n5034);
   registers_reg_5_18_inst : DFF_X1 port map( D => n7553, CK => clk, Q => 
                           n17950, QN => n5035);
   registers_reg_5_17_inst : DFF_X1 port map( D => n7552, CK => clk, Q => 
                           n17949, QN => n5036);
   registers_reg_5_16_inst : DFF_X1 port map( D => n7551, CK => clk, Q => 
                           n17948, QN => n5037);
   registers_reg_5_15_inst : DFF_X1 port map( D => n7550, CK => clk, Q => 
                           n17947, QN => n5038);
   registers_reg_5_14_inst : DFF_X1 port map( D => n7549, CK => clk, Q => 
                           n17946, QN => n5039);
   registers_reg_5_13_inst : DFF_X1 port map( D => n7548, CK => clk, Q => 
                           n17945, QN => n5040);
   registers_reg_5_12_inst : DFF_X1 port map( D => n7547, CK => clk, Q => 
                           n17944, QN => n5041);
   registers_reg_5_11_inst : DFF_X1 port map( D => n7546, CK => clk, Q => 
                           n17943, QN => n5042);
   registers_reg_5_10_inst : DFF_X1 port map( D => n7545, CK => clk, Q => 
                           n17942, QN => n5043);
   registers_reg_5_9_inst : DFF_X1 port map( D => n7544, CK => clk, Q => n17941
                           , QN => n5044);
   registers_reg_5_8_inst : DFF_X1 port map( D => n7543, CK => clk, Q => n17940
                           , QN => n5045);
   registers_reg_5_7_inst : DFF_X1 port map( D => n7542, CK => clk, Q => n17939
                           , QN => n5046);
   registers_reg_5_6_inst : DFF_X1 port map( D => n7541, CK => clk, Q => n17938
                           , QN => n5047);
   registers_reg_5_5_inst : DFF_X1 port map( D => n7540, CK => clk, Q => n17937
                           , QN => n5048);
   registers_reg_5_4_inst : DFF_X1 port map( D => n7539, CK => clk, Q => n17936
                           , QN => n5049);
   registers_reg_6_63_inst : DFF_X1 port map( D => n7662, CK => clk, Q => 
                           n18055, QN => n4924);
   registers_reg_6_62_inst : DFF_X1 port map( D => n7661, CK => clk, Q => 
                           n18054, QN => n4925);
   registers_reg_6_61_inst : DFF_X1 port map( D => n7660, CK => clk, Q => 
                           n18053, QN => n4926);
   registers_reg_6_60_inst : DFF_X1 port map( D => n7659, CK => clk, Q => 
                           n18052, QN => n4927);
   registers_reg_6_59_inst : DFF_X1 port map( D => n7658, CK => clk, Q => 
                           n18051, QN => n4928);
   registers_reg_6_58_inst : DFF_X1 port map( D => n7657, CK => clk, Q => 
                           n18050, QN => n4929);
   registers_reg_6_57_inst : DFF_X1 port map( D => n7656, CK => clk, Q => 
                           n18049, QN => n4930);
   registers_reg_6_56_inst : DFF_X1 port map( D => n7655, CK => clk, Q => 
                           n18048, QN => n4931);
   registers_reg_6_55_inst : DFF_X1 port map( D => n7654, CK => clk, Q => 
                           n18047, QN => n4932);
   registers_reg_6_54_inst : DFF_X1 port map( D => n7653, CK => clk, Q => 
                           n18046, QN => n4933);
   registers_reg_6_53_inst : DFF_X1 port map( D => n7652, CK => clk, Q => 
                           n18045, QN => n4934);
   registers_reg_6_52_inst : DFF_X1 port map( D => n7651, CK => clk, Q => 
                           n18044, QN => n4935);
   registers_reg_6_51_inst : DFF_X1 port map( D => n7650, CK => clk, Q => 
                           n18043, QN => n4936);
   registers_reg_6_50_inst : DFF_X1 port map( D => n7649, CK => clk, Q => 
                           n18042, QN => n4937);
   registers_reg_6_49_inst : DFF_X1 port map( D => n7648, CK => clk, Q => 
                           n18041, QN => n4938);
   registers_reg_6_48_inst : DFF_X1 port map( D => n7647, CK => clk, Q => 
                           n18040, QN => n4939);
   registers_reg_6_47_inst : DFF_X1 port map( D => n7646, CK => clk, Q => 
                           n18039, QN => n4940);
   registers_reg_6_46_inst : DFF_X1 port map( D => n7645, CK => clk, Q => 
                           n18038, QN => n4941);
   registers_reg_6_45_inst : DFF_X1 port map( D => n7644, CK => clk, Q => 
                           n18037, QN => n4942);
   registers_reg_6_44_inst : DFF_X1 port map( D => n7643, CK => clk, Q => 
                           n18036, QN => n4943);
   registers_reg_6_43_inst : DFF_X1 port map( D => n7642, CK => clk, Q => 
                           n18035, QN => n4944);
   registers_reg_6_42_inst : DFF_X1 port map( D => n7641, CK => clk, Q => 
                           n18034, QN => n4945);
   registers_reg_6_41_inst : DFF_X1 port map( D => n7640, CK => clk, Q => 
                           n18033, QN => n4946);
   registers_reg_6_40_inst : DFF_X1 port map( D => n7639, CK => clk, Q => 
                           n18032, QN => n4947);
   registers_reg_6_39_inst : DFF_X1 port map( D => n7638, CK => clk, Q => 
                           n18031, QN => n4948);
   registers_reg_6_38_inst : DFF_X1 port map( D => n7637, CK => clk, Q => 
                           n18030, QN => n4949);
   registers_reg_6_37_inst : DFF_X1 port map( D => n7636, CK => clk, Q => 
                           n18029, QN => n4950);
   registers_reg_6_36_inst : DFF_X1 port map( D => n7635, CK => clk, Q => 
                           n18028, QN => n4951);
   registers_reg_6_35_inst : DFF_X1 port map( D => n7634, CK => clk, Q => 
                           n18027, QN => n4952);
   registers_reg_6_34_inst : DFF_X1 port map( D => n7633, CK => clk, Q => 
                           n18026, QN => n4953);
   registers_reg_6_33_inst : DFF_X1 port map( D => n7632, CK => clk, Q => 
                           n18025, QN => n4954);
   registers_reg_6_32_inst : DFF_X1 port map( D => n7631, CK => clk, Q => 
                           n18024, QN => n4955);
   registers_reg_6_31_inst : DFF_X1 port map( D => n7630, CK => clk, Q => 
                           n18023, QN => n4956);
   registers_reg_6_30_inst : DFF_X1 port map( D => n7629, CK => clk, Q => 
                           n18022, QN => n4957);
   registers_reg_6_29_inst : DFF_X1 port map( D => n7628, CK => clk, Q => 
                           n18021, QN => n4958);
   registers_reg_6_28_inst : DFF_X1 port map( D => n7627, CK => clk, Q => 
                           n18020, QN => n4959);
   registers_reg_6_27_inst : DFF_X1 port map( D => n7626, CK => clk, Q => 
                           n18019, QN => n4960);
   registers_reg_6_26_inst : DFF_X1 port map( D => n7625, CK => clk, Q => 
                           n18018, QN => n4961);
   registers_reg_6_25_inst : DFF_X1 port map( D => n7624, CK => clk, Q => 
                           n18017, QN => n4962);
   registers_reg_6_24_inst : DFF_X1 port map( D => n7623, CK => clk, Q => 
                           n18016, QN => n4963);
   registers_reg_6_23_inst : DFF_X1 port map( D => n7622, CK => clk, Q => 
                           n18015, QN => n4964);
   registers_reg_6_22_inst : DFF_X1 port map( D => n7621, CK => clk, Q => 
                           n18014, QN => n4965);
   registers_reg_6_21_inst : DFF_X1 port map( D => n7620, CK => clk, Q => 
                           n18013, QN => n4966);
   registers_reg_6_20_inst : DFF_X1 port map( D => n7619, CK => clk, Q => 
                           n18012, QN => n4967);
   registers_reg_6_19_inst : DFF_X1 port map( D => n7618, CK => clk, Q => 
                           n18011, QN => n4968);
   registers_reg_6_18_inst : DFF_X1 port map( D => n7617, CK => clk, Q => 
                           n18010, QN => n4969);
   registers_reg_6_17_inst : DFF_X1 port map( D => n7616, CK => clk, Q => 
                           n18009, QN => n4970);
   registers_reg_6_16_inst : DFF_X1 port map( D => n7615, CK => clk, Q => 
                           n18008, QN => n4971);
   registers_reg_6_15_inst : DFF_X1 port map( D => n7614, CK => clk, Q => 
                           n18007, QN => n4972);
   registers_reg_6_14_inst : DFF_X1 port map( D => n7613, CK => clk, Q => 
                           n18006, QN => n4973);
   registers_reg_6_13_inst : DFF_X1 port map( D => n7612, CK => clk, Q => 
                           n18005, QN => n4974);
   registers_reg_6_12_inst : DFF_X1 port map( D => n7611, CK => clk, Q => 
                           n18004, QN => n4975);
   registers_reg_6_11_inst : DFF_X1 port map( D => n7610, CK => clk, Q => 
                           n18003, QN => n4976);
   registers_reg_6_10_inst : DFF_X1 port map( D => n7609, CK => clk, Q => 
                           n18002, QN => n4977);
   registers_reg_6_9_inst : DFF_X1 port map( D => n7608, CK => clk, Q => n18001
                           , QN => n4978);
   registers_reg_6_8_inst : DFF_X1 port map( D => n7607, CK => clk, Q => n18000
                           , QN => n4979);
   registers_reg_6_7_inst : DFF_X1 port map( D => n7606, CK => clk, Q => n17999
                           , QN => n4980);
   registers_reg_6_6_inst : DFF_X1 port map( D => n7605, CK => clk, Q => n17998
                           , QN => n4981);
   registers_reg_6_5_inst : DFF_X1 port map( D => n7604, CK => clk, Q => n17997
                           , QN => n4982);
   registers_reg_6_4_inst : DFF_X1 port map( D => n7603, CK => clk, Q => n17996
                           , QN => n4983);
   registers_reg_20_63_inst : DFF_X1 port map( D => n8558, CK => clk, Q => 
                           n17915, QN => n3974);
   registers_reg_20_62_inst : DFF_X1 port map( D => n8557, CK => clk, Q => 
                           n17914, QN => n3975);
   registers_reg_20_61_inst : DFF_X1 port map( D => n8556, CK => clk, Q => 
                           n17913, QN => n3976);
   registers_reg_20_60_inst : DFF_X1 port map( D => n8555, CK => clk, Q => 
                           n17912, QN => n3977);
   registers_reg_20_59_inst : DFF_X1 port map( D => n8554, CK => clk, Q => 
                           n17887, QN => n3978);
   registers_reg_20_58_inst : DFF_X1 port map( D => n8553, CK => clk, Q => 
                           n17886, QN => n3979);
   registers_reg_20_57_inst : DFF_X1 port map( D => n8552, CK => clk, Q => 
                           n17885, QN => n3980);
   registers_reg_20_56_inst : DFF_X1 port map( D => n8551, CK => clk, Q => 
                           n17884, QN => n3981);
   registers_reg_20_55_inst : DFF_X1 port map( D => n8550, CK => clk, Q => 
                           n17883, QN => n3982);
   registers_reg_20_54_inst : DFF_X1 port map( D => n8549, CK => clk, Q => 
                           n17882, QN => n3983);
   registers_reg_20_53_inst : DFF_X1 port map( D => n8548, CK => clk, Q => 
                           n17881, QN => n3984);
   registers_reg_20_52_inst : DFF_X1 port map( D => n8547, CK => clk, Q => 
                           n17880, QN => n3985);
   registers_reg_20_51_inst : DFF_X1 port map( D => n8546, CK => clk, Q => 
                           n17879, QN => n3986);
   registers_reg_20_50_inst : DFF_X1 port map( D => n8545, CK => clk, Q => 
                           n17878, QN => n3987);
   registers_reg_20_49_inst : DFF_X1 port map( D => n8544, CK => clk, Q => 
                           n17877, QN => n3988);
   registers_reg_20_48_inst : DFF_X1 port map( D => n8543, CK => clk, Q => 
                           n17876, QN => n3989);
   registers_reg_20_47_inst : DFF_X1 port map( D => n8542, CK => clk, Q => 
                           n17924, QN => n3990);
   registers_reg_20_46_inst : DFF_X1 port map( D => n8541, CK => clk, Q => 
                           n17923, QN => n3991);
   registers_reg_20_45_inst : DFF_X1 port map( D => n8540, CK => clk, Q => 
                           n17922, QN => n3992);
   registers_reg_20_44_inst : DFF_X1 port map( D => n8539, CK => clk, Q => 
                           n17921, QN => n3993);
   registers_reg_20_43_inst : DFF_X1 port map( D => n8538, CK => clk, Q => 
                           n17920, QN => n3994);
   registers_reg_20_42_inst : DFF_X1 port map( D => n8537, CK => clk, Q => 
                           n17919, QN => n3995);
   registers_reg_20_41_inst : DFF_X1 port map( D => n8536, CK => clk, Q => 
                           n17918, QN => n3996);
   registers_reg_20_40_inst : DFF_X1 port map( D => n8535, CK => clk, Q => 
                           n17917, QN => n3997);
   registers_reg_20_39_inst : DFF_X1 port map( D => n8534, CK => clk, Q => 
                           n17916, QN => n3998);
   registers_reg_20_38_inst : DFF_X1 port map( D => n8533, CK => clk, Q => 
                           n17935, QN => n3999);
   registers_reg_20_37_inst : DFF_X1 port map( D => n8532, CK => clk, Q => 
                           n17926, QN => n4000);
   registers_reg_20_36_inst : DFF_X1 port map( D => n8531, CK => clk, Q => 
                           n17925, QN => n4001);
   registers_reg_20_35_inst : DFF_X1 port map( D => n8530, CK => clk, Q => 
                           n17911, QN => n4002);
   registers_reg_20_34_inst : DFF_X1 port map( D => n8529, CK => clk, Q => 
                           n17910, QN => n4003);
   registers_reg_20_33_inst : DFF_X1 port map( D => n8528, CK => clk, Q => 
                           n17909, QN => n4004);
   registers_reg_20_32_inst : DFF_X1 port map( D => n8527, CK => clk, Q => 
                           n17908, QN => n4005);
   registers_reg_20_31_inst : DFF_X1 port map( D => n8526, CK => clk, Q => 
                           n17907, QN => n4006);
   registers_reg_20_30_inst : DFF_X1 port map( D => n8525, CK => clk, Q => 
                           n17906, QN => n4007);
   registers_reg_20_29_inst : DFF_X1 port map( D => n8524, CK => clk, Q => 
                           n17905, QN => n4008);
   registers_reg_20_28_inst : DFF_X1 port map( D => n8523, CK => clk, Q => 
                           n17904, QN => n4009);
   registers_reg_20_27_inst : DFF_X1 port map( D => n8522, CK => clk, Q => 
                           n17903, QN => n4010);
   registers_reg_20_26_inst : DFF_X1 port map( D => n8521, CK => clk, Q => 
                           n17902, QN => n4011);
   registers_reg_20_25_inst : DFF_X1 port map( D => n8520, CK => clk, Q => 
                           n17901, QN => n4012);
   registers_reg_20_24_inst : DFF_X1 port map( D => n8519, CK => clk, Q => 
                           n17900, QN => n4013);
   registers_reg_20_23_inst : DFF_X1 port map( D => n8518, CK => clk, Q => 
                           n17899, QN => n4014);
   registers_reg_20_22_inst : DFF_X1 port map( D => n8517, CK => clk, Q => 
                           n17898, QN => n4015);
   registers_reg_20_21_inst : DFF_X1 port map( D => n8516, CK => clk, Q => 
                           n17897, QN => n4016);
   registers_reg_20_20_inst : DFF_X1 port map( D => n8515, CK => clk, Q => 
                           n17896, QN => n4017);
   registers_reg_20_19_inst : DFF_X1 port map( D => n8514, CK => clk, Q => 
                           n17895, QN => n4018);
   registers_reg_20_18_inst : DFF_X1 port map( D => n8513, CK => clk, Q => 
                           n17894, QN => n4019);
   registers_reg_20_17_inst : DFF_X1 port map( D => n8512, CK => clk, Q => 
                           n17893, QN => n4020);
   registers_reg_20_16_inst : DFF_X1 port map( D => n8511, CK => clk, Q => 
                           n17892, QN => n4021);
   registers_reg_20_15_inst : DFF_X1 port map( D => n8510, CK => clk, Q => 
                           n17891, QN => n4022);
   registers_reg_20_14_inst : DFF_X1 port map( D => n8509, CK => clk, Q => 
                           n17890, QN => n4023);
   registers_reg_20_13_inst : DFF_X1 port map( D => n8508, CK => clk, Q => 
                           n17889, QN => n4024);
   registers_reg_20_12_inst : DFF_X1 port map( D => n8507, CK => clk, Q => 
                           n17888, QN => n4025);
   registers_reg_20_11_inst : DFF_X1 port map( D => n8506, CK => clk, Q => 
                           n17934, QN => n4026);
   registers_reg_20_10_inst : DFF_X1 port map( D => n8505, CK => clk, Q => 
                           n17933, QN => n4027);
   registers_reg_20_9_inst : DFF_X1 port map( D => n8504, CK => clk, Q => 
                           n17932, QN => n4028);
   registers_reg_20_8_inst : DFF_X1 port map( D => n8503, CK => clk, Q => 
                           n17931, QN => n4029);
   registers_reg_20_7_inst : DFF_X1 port map( D => n8502, CK => clk, Q => 
                           n17930, QN => n4030);
   registers_reg_20_6_inst : DFF_X1 port map( D => n8501, CK => clk, Q => 
                           n17929, QN => n4031);
   registers_reg_20_5_inst : DFF_X1 port map( D => n8500, CK => clk, Q => 
                           n17928, QN => n4032);
   registers_reg_20_4_inst : DFF_X1 port map( D => n8499, CK => clk, Q => 
                           n17927, QN => n4033);
   registers_reg_23_63_inst : DFF_X1 port map( D => n8750, CK => clk, Q => 
                           n_1066, QN => n3773);
   registers_reg_23_62_inst : DFF_X1 port map( D => n8749, CK => clk, Q => 
                           n_1067, QN => n3774);
   registers_reg_23_61_inst : DFF_X1 port map( D => n8748, CK => clk, Q => 
                           n_1068, QN => n3775);
   registers_reg_23_60_inst : DFF_X1 port map( D => n8747, CK => clk, Q => 
                           n_1069, QN => n3776);
   registers_reg_23_59_inst : DFF_X1 port map( D => n8746, CK => clk, Q => 
                           n_1070, QN => n3777);
   registers_reg_23_58_inst : DFF_X1 port map( D => n8745, CK => clk, Q => 
                           n_1071, QN => n3778);
   registers_reg_23_57_inst : DFF_X1 port map( D => n8744, CK => clk, Q => 
                           n_1072, QN => n3779);
   registers_reg_23_56_inst : DFF_X1 port map( D => n8743, CK => clk, Q => 
                           n_1073, QN => n3780);
   registers_reg_23_55_inst : DFF_X1 port map( D => n8742, CK => clk, Q => 
                           n_1074, QN => n3781);
   registers_reg_23_54_inst : DFF_X1 port map( D => n8741, CK => clk, Q => 
                           n_1075, QN => n3782);
   registers_reg_23_53_inst : DFF_X1 port map( D => n8740, CK => clk, Q => 
                           n_1076, QN => n3783);
   registers_reg_23_52_inst : DFF_X1 port map( D => n8739, CK => clk, Q => 
                           n_1077, QN => n3784);
   registers_reg_23_51_inst : DFF_X1 port map( D => n8738, CK => clk, Q => 
                           n_1078, QN => n3785);
   registers_reg_23_50_inst : DFF_X1 port map( D => n8737, CK => clk, Q => 
                           n_1079, QN => n3786);
   registers_reg_23_49_inst : DFF_X1 port map( D => n8736, CK => clk, Q => 
                           n_1080, QN => n3787);
   registers_reg_23_48_inst : DFF_X1 port map( D => n8735, CK => clk, Q => 
                           n_1081, QN => n3788);
   registers_reg_23_47_inst : DFF_X1 port map( D => n8734, CK => clk, Q => 
                           n_1082, QN => n3789);
   registers_reg_23_46_inst : DFF_X1 port map( D => n8733, CK => clk, Q => 
                           n_1083, QN => n3790);
   registers_reg_23_45_inst : DFF_X1 port map( D => n8732, CK => clk, Q => 
                           n_1084, QN => n3791);
   registers_reg_23_44_inst : DFF_X1 port map( D => n8731, CK => clk, Q => 
                           n_1085, QN => n3792);
   registers_reg_23_43_inst : DFF_X1 port map( D => n8730, CK => clk, Q => 
                           n_1086, QN => n3793);
   registers_reg_23_42_inst : DFF_X1 port map( D => n8729, CK => clk, Q => 
                           n_1087, QN => n3794);
   registers_reg_23_41_inst : DFF_X1 port map( D => n8728, CK => clk, Q => 
                           n_1088, QN => n3795);
   registers_reg_23_40_inst : DFF_X1 port map( D => n8727, CK => clk, Q => 
                           n_1089, QN => n3796);
   registers_reg_23_39_inst : DFF_X1 port map( D => n8726, CK => clk, Q => 
                           n_1090, QN => n3797);
   registers_reg_23_38_inst : DFF_X1 port map( D => n8725, CK => clk, Q => 
                           n_1091, QN => n3798);
   registers_reg_23_37_inst : DFF_X1 port map( D => n8724, CK => clk, Q => 
                           n_1092, QN => n3799);
   registers_reg_23_36_inst : DFF_X1 port map( D => n8723, CK => clk, Q => 
                           n_1093, QN => n3800);
   registers_reg_23_35_inst : DFF_X1 port map( D => n8722, CK => clk, Q => 
                           n_1094, QN => n3801);
   registers_reg_23_34_inst : DFF_X1 port map( D => n8721, CK => clk, Q => 
                           n_1095, QN => n3802);
   registers_reg_23_33_inst : DFF_X1 port map( D => n8720, CK => clk, Q => 
                           n_1096, QN => n3803);
   registers_reg_23_32_inst : DFF_X1 port map( D => n8719, CK => clk, Q => 
                           n_1097, QN => n3804);
   registers_reg_23_31_inst : DFF_X1 port map( D => n8718, CK => clk, Q => 
                           n_1098, QN => n3805);
   registers_reg_23_30_inst : DFF_X1 port map( D => n8717, CK => clk, Q => 
                           n_1099, QN => n3806);
   registers_reg_23_29_inst : DFF_X1 port map( D => n8716, CK => clk, Q => 
                           n_1100, QN => n3807);
   registers_reg_23_28_inst : DFF_X1 port map( D => n8715, CK => clk, Q => 
                           n_1101, QN => n3808);
   registers_reg_23_27_inst : DFF_X1 port map( D => n8714, CK => clk, Q => 
                           n_1102, QN => n3809);
   registers_reg_23_26_inst : DFF_X1 port map( D => n8713, CK => clk, Q => 
                           n_1103, QN => n3810);
   registers_reg_23_25_inst : DFF_X1 port map( D => n8712, CK => clk, Q => 
                           n_1104, QN => n3811);
   registers_reg_23_24_inst : DFF_X1 port map( D => n8711, CK => clk, Q => 
                           n_1105, QN => n3812);
   registers_reg_23_23_inst : DFF_X1 port map( D => n8710, CK => clk, Q => 
                           n_1106, QN => n3813);
   registers_reg_23_22_inst : DFF_X1 port map( D => n8709, CK => clk, Q => 
                           n_1107, QN => n3814);
   registers_reg_23_21_inst : DFF_X1 port map( D => n8708, CK => clk, Q => 
                           n_1108, QN => n3815);
   registers_reg_23_20_inst : DFF_X1 port map( D => n8707, CK => clk, Q => 
                           n_1109, QN => n3816);
   registers_reg_23_19_inst : DFF_X1 port map( D => n8706, CK => clk, Q => 
                           n_1110, QN => n3817);
   registers_reg_23_18_inst : DFF_X1 port map( D => n8705, CK => clk, Q => 
                           n_1111, QN => n3818);
   registers_reg_23_17_inst : DFF_X1 port map( D => n8704, CK => clk, Q => 
                           n_1112, QN => n3819);
   registers_reg_23_16_inst : DFF_X1 port map( D => n8703, CK => clk, Q => 
                           n_1113, QN => n3820);
   registers_reg_23_15_inst : DFF_X1 port map( D => n8702, CK => clk, Q => 
                           n_1114, QN => n3821);
   registers_reg_23_14_inst : DFF_X1 port map( D => n8701, CK => clk, Q => 
                           n_1115, QN => n3822);
   registers_reg_23_13_inst : DFF_X1 port map( D => n8700, CK => clk, Q => 
                           n_1116, QN => n3823);
   registers_reg_23_12_inst : DFF_X1 port map( D => n8699, CK => clk, Q => 
                           n_1117, QN => n3824);
   registers_reg_23_11_inst : DFF_X1 port map( D => n8698, CK => clk, Q => 
                           n_1118, QN => n3825);
   registers_reg_23_10_inst : DFF_X1 port map( D => n8697, CK => clk, Q => 
                           n_1119, QN => n3826);
   registers_reg_23_9_inst : DFF_X1 port map( D => n8696, CK => clk, Q => 
                           n_1120, QN => n3827);
   registers_reg_23_8_inst : DFF_X1 port map( D => n8695, CK => clk, Q => 
                           n_1121, QN => n3828);
   registers_reg_23_7_inst : DFF_X1 port map( D => n8694, CK => clk, Q => 
                           n_1122, QN => n3829);
   registers_reg_23_6_inst : DFF_X1 port map( D => n8693, CK => clk, Q => 
                           n_1123, QN => n3830);
   registers_reg_23_5_inst : DFF_X1 port map( D => n8692, CK => clk, Q => 
                           n_1124, QN => n3831);
   registers_reg_23_4_inst : DFF_X1 port map( D => n8691, CK => clk, Q => 
                           n_1125, QN => n3832);
   out_to_mem_reg_2_inst : DFF_X1 port map( D => n7031, CK => clk, Q => 
                           out_to_mem_2_port, QN => n15079);
   out_to_mem_reg_1_inst : DFF_X1 port map( D => n7027, CK => clk, Q => 
                           out_to_mem_1_port, QN => n15078);
   out_to_mem_reg_0_inst : DFF_X1 port map( D => n7023, CK => clk, Q => 
                           out_to_mem_0_port, QN => n15077);
   registers_reg_7_63_inst : DFF_X1 port map( D => n7726, CK => clk, Q => 
                           n18179, QN => n4858);
   registers_reg_7_62_inst : DFF_X1 port map( D => n7725, CK => clk, Q => 
                           n18178, QN => n4859);
   registers_reg_7_61_inst : DFF_X1 port map( D => n7724, CK => clk, Q => 
                           n18177, QN => n4860);
   registers_reg_7_60_inst : DFF_X1 port map( D => n7723, CK => clk, Q => 
                           n18176, QN => n4861);
   registers_reg_7_59_inst : DFF_X1 port map( D => n7722, CK => clk, Q => 
                           n18201, QN => n4862);
   registers_reg_7_58_inst : DFF_X1 port map( D => n7721, CK => clk, Q => 
                           n18200, QN => n4863);
   registers_reg_7_57_inst : DFF_X1 port map( D => n7720, CK => clk, Q => 
                           n18199, QN => n4864);
   registers_reg_7_56_inst : DFF_X1 port map( D => n7719, CK => clk, Q => 
                           n18198, QN => n4865);
   registers_reg_7_55_inst : DFF_X1 port map( D => n7718, CK => clk, Q => 
                           n18197, QN => n4866);
   registers_reg_7_54_inst : DFF_X1 port map( D => n7717, CK => clk, Q => 
                           n18196, QN => n4867);
   registers_reg_7_53_inst : DFF_X1 port map( D => n7716, CK => clk, Q => 
                           n18195, QN => n4868);
   registers_reg_7_52_inst : DFF_X1 port map( D => n7715, CK => clk, Q => 
                           n18194, QN => n4869);
   registers_reg_7_51_inst : DFF_X1 port map( D => n7714, CK => clk, Q => 
                           n18193, QN => n4870);
   registers_reg_7_50_inst : DFF_X1 port map( D => n7713, CK => clk, Q => 
                           n18192, QN => n4871);
   registers_reg_7_49_inst : DFF_X1 port map( D => n7712, CK => clk, Q => 
                           n18191, QN => n4872);
   registers_reg_7_48_inst : DFF_X1 port map( D => n7711, CK => clk, Q => 
                           n18190, QN => n4873);
   registers_reg_7_47_inst : DFF_X1 port map( D => n7710, CK => clk, Q => 
                           n18189, QN => n4874);
   registers_reg_7_46_inst : DFF_X1 port map( D => n7709, CK => clk, Q => 
                           n18188, QN => n4875);
   registers_reg_7_45_inst : DFF_X1 port map( D => n7708, CK => clk, Q => 
                           n18187, QN => n4876);
   registers_reg_7_44_inst : DFF_X1 port map( D => n7707, CK => clk, Q => 
                           n18186, QN => n4877);
   registers_reg_7_43_inst : DFF_X1 port map( D => n7706, CK => clk, Q => 
                           n18185, QN => n4878);
   registers_reg_7_42_inst : DFF_X1 port map( D => n7705, CK => clk, Q => 
                           n18184, QN => n4879);
   registers_reg_7_41_inst : DFF_X1 port map( D => n7704, CK => clk, Q => 
                           n18183, QN => n4880);
   registers_reg_7_40_inst : DFF_X1 port map( D => n7703, CK => clk, Q => 
                           n18182, QN => n4881);
   registers_reg_7_39_inst : DFF_X1 port map( D => n7702, CK => clk, Q => 
                           n18181, QN => n4882);
   registers_reg_7_38_inst : DFF_X1 port map( D => n7701, CK => clk, Q => 
                           n18180, QN => n4883);
   registers_reg_7_37_inst : DFF_X1 port map( D => n7700, CK => clk, Q => 
                           n18235, QN => n4884);
   registers_reg_7_36_inst : DFF_X1 port map( D => n7699, CK => clk, Q => 
                           n18234, QN => n4885);
   registers_reg_7_35_inst : DFF_X1 port map( D => n7698, CK => clk, Q => 
                           n18233, QN => n4886);
   registers_reg_7_34_inst : DFF_X1 port map( D => n7697, CK => clk, Q => 
                           n18232, QN => n4887);
   registers_reg_7_33_inst : DFF_X1 port map( D => n7696, CK => clk, Q => 
                           n18231, QN => n4888);
   registers_reg_7_32_inst : DFF_X1 port map( D => n7695, CK => clk, Q => 
                           n18230, QN => n4889);
   registers_reg_7_31_inst : DFF_X1 port map( D => n7694, CK => clk, Q => 
                           n18229, QN => n4890);
   registers_reg_7_30_inst : DFF_X1 port map( D => n7693, CK => clk, Q => 
                           n18228, QN => n4891);
   registers_reg_7_29_inst : DFF_X1 port map( D => n7692, CK => clk, Q => 
                           n18227, QN => n4892);
   registers_reg_7_28_inst : DFF_X1 port map( D => n7691, CK => clk, Q => 
                           n18226, QN => n4893);
   registers_reg_7_27_inst : DFF_X1 port map( D => n7690, CK => clk, Q => 
                           n18225, QN => n4894);
   registers_reg_7_26_inst : DFF_X1 port map( D => n7689, CK => clk, Q => 
                           n18224, QN => n4895);
   registers_reg_7_25_inst : DFF_X1 port map( D => n7688, CK => clk, Q => 
                           n18223, QN => n4896);
   registers_reg_7_24_inst : DFF_X1 port map( D => n7687, CK => clk, Q => 
                           n18222, QN => n4897);
   registers_reg_7_23_inst : DFF_X1 port map( D => n7686, CK => clk, Q => 
                           n18221, QN => n4898);
   registers_reg_7_22_inst : DFF_X1 port map( D => n7685, CK => clk, Q => 
                           n18220, QN => n4899);
   registers_reg_7_21_inst : DFF_X1 port map( D => n7684, CK => clk, Q => 
                           n18219, QN => n4900);
   registers_reg_7_20_inst : DFF_X1 port map( D => n7683, CK => clk, Q => 
                           n18218, QN => n4901);
   registers_reg_7_19_inst : DFF_X1 port map( D => n7682, CK => clk, Q => 
                           n18217, QN => n4902);
   registers_reg_7_18_inst : DFF_X1 port map( D => n7681, CK => clk, Q => 
                           n18216, QN => n4903);
   registers_reg_7_17_inst : DFF_X1 port map( D => n7680, CK => clk, Q => 
                           n18215, QN => n4904);
   registers_reg_7_16_inst : DFF_X1 port map( D => n7679, CK => clk, Q => 
                           n18214, QN => n4905);
   registers_reg_7_15_inst : DFF_X1 port map( D => n7678, CK => clk, Q => 
                           n18213, QN => n4906);
   registers_reg_7_14_inst : DFF_X1 port map( D => n7677, CK => clk, Q => 
                           n18212, QN => n4907);
   registers_reg_7_13_inst : DFF_X1 port map( D => n7676, CK => clk, Q => 
                           n18211, QN => n4908);
   registers_reg_7_12_inst : DFF_X1 port map( D => n7675, CK => clk, Q => 
                           n18210, QN => n4909);
   registers_reg_7_11_inst : DFF_X1 port map( D => n7674, CK => clk, Q => 
                           n18209, QN => n4910);
   registers_reg_7_10_inst : DFF_X1 port map( D => n7673, CK => clk, Q => 
                           n18208, QN => n4911);
   registers_reg_7_9_inst : DFF_X1 port map( D => n7672, CK => clk, Q => n18207
                           , QN => n4912);
   registers_reg_7_8_inst : DFF_X1 port map( D => n7671, CK => clk, Q => n18206
                           , QN => n4913);
   registers_reg_7_7_inst : DFF_X1 port map( D => n7670, CK => clk, Q => n18205
                           , QN => n4914);
   registers_reg_7_6_inst : DFF_X1 port map( D => n7669, CK => clk, Q => n18204
                           , QN => n4915);
   registers_reg_7_5_inst : DFF_X1 port map( D => n7668, CK => clk, Q => n18203
                           , QN => n4916);
   registers_reg_7_4_inst : DFF_X1 port map( D => n7667, CK => clk, Q => n18202
                           , QN => n4917);
   n4 <= '0';
   n5 <= '0';
   n6 <= '0';
   U1725 : NAND2_X2 port map( A1 => n2216, A2 => n2219, ZN => n1715);
   U2055 : OR2_X2 port map( A1 => n2375, A2 => n2092, ZN => n1726);
   U7374 : INV_X2 port map( A => n11702, ZN => n11681);
   U7403 : AOI21_X2 port map( B1 => n11751, B2 => sub_123_carry_4_port, A => 
                           n11748, ZN => n1940);
   U7439 : NAND3_X1 port map( A1 => n1870, A2 => n1871, A3 => count3(0), ZN => 
                           n1697);
   U7440 : NAND3_X1 port map( A1 => n1871, A2 => n1939, A3 => n1870, ZN => 
                           n1705);
   U7441 : NAND3_X1 port map( A1 => n1870, A2 => count3(0), A3 => n1943, ZN => 
                           n1708);
   U7442 : NAND3_X1 port map( A1 => n1870, A2 => n1939, A3 => n1943, ZN => 
                           n1712);
   U7443 : NAND3_X1 port map( A1 => N148, A2 => N150, A3 => n2087, ZN => n1700)
                           ;
   U7444 : NAND3_X1 port map( A1 => N150, A2 => n2094, A3 => n2087, ZN => n1704
                           );
   U7445 : NAND3_X1 port map( A1 => N148, A2 => n2207, A3 => n2087, ZN => n1716
                           );
   U7446 : NAND3_X1 port map( A1 => n2094, A2 => n2207, A3 => n2087, ZN => 
                           n1719);
   U7447 : NAND3_X1 port map( A1 => N148, A2 => N150, A3 => n2252, ZN => n1727)
                           ;
   U7448 : NAND3_X1 port map( A1 => N150, A2 => n2094, A3 => n2252, ZN => n1797
                           );
   U7449 : NAND3_X1 port map( A1 => N148, A2 => n2207, A3 => n2252, ZN => n1869
                           );
   U7450 : NAND3_X1 port map( A1 => n2093, A2 => n2219, A3 => n2091, ZN => 
                           n1868);
   U7451 : NAND3_X1 port map( A1 => n2094, A2 => n2207, A3 => n2252, ZN => 
                           n1938);
   U7452 : NAND3_X1 port map( A1 => n11673, A2 => n11674, A3 => n11675, ZN => 
                           n3148);
   U7453 : NAND3_X1 port map( A1 => n11680, A2 => n11683, A3 => n11675, ZN => 
                           n3172);
   U7454 : NAND3_X1 port map( A1 => n11675, A2 => n11674, A3 => n11700, ZN => 
                           n3170);
   U7455 : NAND3_X1 port map( A1 => n1946, A2 => n1939, A3 => n1871, ZN => 
                           n2082);
   U7456 : NAND3_X1 port map( A1 => n1946, A2 => n1939, A3 => n1943, ZN => 
                           n2090);
   U7457 : NAND3_X1 port map( A1 => n11680, A2 => n2093, A3 => n11718, ZN => 
                           n11696);
   U7458 : NAND3_X1 port map( A1 => n11680, A2 => n11716, A3 => n11718, ZN => 
                           n11710);
   U7460 : NAND3_X1 port map( A1 => n11674, A2 => n2093, A3 => n11718, ZN => 
                           n11708);
   U7461 : NAND3_X1 port map( A1 => n2091, A2 => n2093, A3 => n18902, ZN => 
                           n11694);
   U7462 : XOR2_X1 port map( A => n11722, B => n11723, Z => n2091);
   U7463 : NAND3_X1 port map( A1 => n1871, A2 => n1946, A3 => count3(0), ZN => 
                           n2015);
   U7465 : XOR2_X1 port map( A => n11743, B => n11739, Z => n11671);
   U7466 : NAND3_X1 port map( A1 => n11716, A2 => n11674, A3 => n11718, ZN => 
                           n11686);
   U7467 : XOR2_X1 port map( A => count3(1), B => n11753, Z => n11680);
   U7468 : XOR2_X1 port map( A => n11732, B => n11755, Z => n2093);
   r507 : register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_2 port map( A(4) 
                           => add_rd2(4), A(3) => add_rd2(3), A(2) => 
                           add_rd2(2), A(1) => add_rd2(1), A(0) => add_rd2(0), 
                           B(4) => U3_U4_Z_4, B(3) => U3_U4_Z_3, B(2) => 
                           U3_U4_Z_2, B(1) => U3_U4_Z_1, B(0) => U3_U4_Z_0, CI 
                           => n4, SUM(4) => N127, SUM(3) => 
                           sub_105_carry_4_port, SUM(2) => N115, SUM(1) => N114
                           , SUM(0) => N113, CO => n1748);
   r497 : register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_3 port map( A(4) 
                           => add_rd1(4), A(3) => add_rd1(3), A(2) => 
                           add_rd1(2), A(1) => add_rd1(1), A(0) => add_rd1(0), 
                           B(4) => U3_U2_Z_4, B(3) => U3_U2_Z_3, B(2) => 
                           U3_U2_Z_2, B(1) => U3_U2_Z_1, B(0) => U3_U2_Z_0, CI 
                           => n5, SUM(4) => N92, SUM(3) => sub_86_carry_4_port,
                           SUM(2) => N80, SUM(1) => N79, SUM(0) => N78, CO => 
                           n1747);
   r517 : register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_add_4 port map( A(4) 
                           => add_wr(4), A(3) => add_wr(3), A(2) => add_wr(2), 
                           A(1) => add_wr(1), A(0) => add_wr(0), B(4) => 
                           U3_U6_Z_4, B(3) => U3_U6_Z_3, B(2) => U3_U6_Z_2, 
                           B(1) => U3_U6_Z_1, B(0) => U3_U6_Z_0, CI => n6, 
                           SUM(4) => N162, SUM(3) => sub_123_carry_4_port, 
                           SUM(2) => N150, SUM(1) => N149, SUM(0) => N148, CO 
                           => n1746);
   registers_reg_13_3_inst : DFF_X1 port map( D => n8050, CK => clk, Q => 
                           n11416, QN => n4508);
   registers_reg_13_2_inst : DFF_X1 port map( D => n8049, CK => clk, Q => 
                           n11483, QN => n4509);
   registers_reg_13_1_inst : DFF_X1 port map( D => n8048, CK => clk, Q => 
                           n11551, QN => n4510);
   registers_reg_13_0_inst : DFF_X1 port map( D => n8047, CK => clk, Q => 
                           n11712, QN => n4511);
   registers_reg_12_3_inst : DFF_X1 port map( D => n7986, CK => clk, Q => 
                           n18901, QN => n4577);
   registers_reg_12_2_inst : DFF_X1 port map( D => n7985, CK => clk, Q => 
                           n18900, QN => n4578);
   registers_reg_12_1_inst : DFF_X1 port map( D => n7984, CK => clk, Q => 
                           n18899, QN => n4579);
   registers_reg_12_0_inst : DFF_X1 port map( D => n7983, CK => clk, Q => 
                           n18898, QN => n4580);
   registers_reg_10_3_inst : DFF_X1 port map( D => n7858, CK => clk, Q => 
                           n11411, QN => n4714);
   registers_reg_10_2_inst : DFF_X1 port map( D => n7857, CK => clk, Q => 
                           n11478, QN => n4715);
   registers_reg_10_1_inst : DFF_X1 port map( D => n7856, CK => clk, Q => 
                           n11546, QN => n4716);
   registers_reg_9_3_inst : DFF_X1 port map( D => n7794, CK => clk, Q => n11379
                           , QN => n4780);
   registers_reg_9_2_inst : DFF_X1 port map( D => n7793, CK => clk, Q => n11447
                           , QN => n4781);
   registers_reg_9_1_inst : DFF_X1 port map( D => n7792, CK => clk, Q => n11514
                           , QN => n4782);
   registers_reg_8_3_inst : DFF_X1 port map( D => n7730, CK => clk, Q => n11417
                           , QN => n4847);
   registers_reg_8_2_inst : DFF_X1 port map( D => n7729, CK => clk, Q => n11484
                           , QN => n4848);
   registers_reg_8_1_inst : DFF_X1 port map( D => n7728, CK => clk, Q => n11552
                           , QN => n4849);
   registers_reg_10_0_inst : DFF_X1 port map( D => n7855, CK => clk, Q => 
                           n11690, QN => n4717);
   registers_reg_9_0_inst : DFF_X1 port map( D => n7791, CK => clk, Q => n11619
                           , QN => n4783);
   registers_reg_8_0_inst : DFF_X1 port map( D => n7727, CK => clk, Q => n11713
                           , QN => n4850);
   registers_reg_1_3_inst : DFF_X1 port map( D => n7282, CK => clk, Q => n18897
                           , QN => n5901);
   registers_reg_1_2_inst : DFF_X1 port map( D => n7281, CK => clk, Q => n18896
                           , QN => n5966);
   registers_reg_1_1_inst : DFF_X1 port map( D => n7280, CK => clk, Q => n18895
                           , QN => n5968);
   registers_reg_1_0_inst : DFF_X1 port map( D => n7279, CK => clk, Q => n18894
                           , QN => n6033);
   registers_reg_24_3_inst : DFF_X1 port map( D => n8754, CK => clk, Q => 
                           n11368, QN => n3767);
   registers_reg_24_2_inst : DFF_X1 port map( D => n8753, CK => clk, Q => 
                           n11435, QN => n3768);
   registers_reg_24_1_inst : DFF_X1 port map( D => n8752, CK => clk, Q => 
                           n11503, QN => n3769);
   registers_reg_24_0_inst : DFF_X1 port map( D => n8751, CK => clk, Q => 
                           n11598, QN => n3770);
   registers_reg_16_3_inst : DFF_X1 port map( D => n8242, CK => clk, Q => 
                           n11378, QN => n4306);
   registers_reg_16_2_inst : DFF_X1 port map( D => n8241, CK => clk, Q => 
                           n11446, QN => n4307);
   registers_reg_16_1_inst : DFF_X1 port map( D => n8240, CK => clk, Q => 
                           n11513, QN => n4308);
   registers_reg_16_0_inst : DFF_X1 port map( D => n8239, CK => clk, Q => 
                           n11618, QN => n4309);
   registers_reg_28_3_inst : DFF_X1 port map( D => n9010, CK => clk, Q => 
                           n18893, QN => n3499);
   registers_reg_28_2_inst : DFF_X1 port map( D => n9009, CK => clk, Q => 
                           n18892, QN => n3500);
   registers_reg_28_1_inst : DFF_X1 port map( D => n9008, CK => clk, Q => 
                           n18891, QN => n3501);
   registers_reg_28_0_inst : DFF_X1 port map( D => n9007, CK => clk, Q => 
                           n18890, QN => n3502);
   registers_reg_26_3_inst : DFF_X1 port map( D => n8882, CK => clk, Q => 
                           n18889, QN => n3634);
   registers_reg_26_2_inst : DFF_X1 port map( D => n8881, CK => clk, Q => 
                           n18888, QN => n3635);
   registers_reg_26_1_inst : DFF_X1 port map( D => n8880, CK => clk, Q => 
                           n18887, QN => n3636);
   registers_reg_26_0_inst : DFF_X1 port map( D => n8879, CK => clk, Q => 
                           n18886, QN => n3637);
   registers_reg_13_63_inst : DFF_X1 port map( D => n8110, CK => clk, Q => 
                           n3188, QN => n4448);
   registers_reg_13_62_inst : DFF_X1 port map( D => n8109, CK => clk, Q => 
                           n3570, QN => n4449);
   registers_reg_13_61_inst : DFF_X1 port map( D => n8108, CK => clk, Q => 
                           n4852, QN => n4450);
   registers_reg_13_60_inst : DFF_X1 port map( D => n8107, CK => clk, Q => 
                           n5337, QN => n4451);
   registers_reg_13_59_inst : DFF_X1 port map( D => n8106, CK => clk, Q => 
                           n5407, QN => n4452);
   registers_reg_13_58_inst : DFF_X1 port map( D => n8105, CK => clk, Q => 
                           n5475, QN => n4453);
   registers_reg_13_57_inst : DFF_X1 port map( D => n8104, CK => clk, Q => 
                           n5544, QN => n4454);
   registers_reg_13_56_inst : DFF_X1 port map( D => n8103, CK => clk, Q => 
                           n5613, QN => n4455);
   registers_reg_13_55_inst : DFF_X1 port map( D => n8102, CK => clk, Q => 
                           n5681, QN => n4456);
   registers_reg_13_54_inst : DFF_X1 port map( D => n8101, CK => clk, Q => 
                           n5751, QN => n4457);
   registers_reg_13_53_inst : DFF_X1 port map( D => n8100, CK => clk, Q => 
                           n5823, QN => n4458);
   registers_reg_13_52_inst : DFF_X1 port map( D => n8099, CK => clk, Q => 
                           n5890, QN => n4459);
   registers_reg_13_51_inst : DFF_X1 port map( D => n8098, CK => clk, Q => 
                           n5957, QN => n4460);
   registers_reg_13_50_inst : DFF_X1 port map( D => n8097, CK => clk, Q => 
                           n6025, QN => n4461);
   registers_reg_13_49_inst : DFF_X1 port map( D => n8096, CK => clk, Q => 
                           n6093, QN => n4462);
   registers_reg_13_48_inst : DFF_X1 port map( D => n8095, CK => clk, Q => 
                           n6159, QN => n4463);
   registers_reg_13_47_inst : DFF_X1 port map( D => n8094, CK => clk, Q => 
                           n6225, QN => n4464);
   registers_reg_13_46_inst : DFF_X1 port map( D => n8093, CK => clk, Q => 
                           n6291, QN => n4465);
   registers_reg_13_45_inst : DFF_X1 port map( D => n8092, CK => clk, Q => 
                           n6357, QN => n4466);
   registers_reg_13_44_inst : DFF_X1 port map( D => n8091, CK => clk, Q => 
                           n6423, QN => n4467);
   registers_reg_13_43_inst : DFF_X1 port map( D => n8090, CK => clk, Q => 
                           n6489, QN => n4468);
   registers_reg_13_42_inst : DFF_X1 port map( D => n8089, CK => clk, Q => 
                           n6555, QN => n4469);
   registers_reg_13_41_inst : DFF_X1 port map( D => n8088, CK => clk, Q => 
                           n6621, QN => n4470);
   registers_reg_13_40_inst : DFF_X1 port map( D => n8087, CK => clk, Q => 
                           n6688, QN => n4471);
   registers_reg_13_39_inst : DFF_X1 port map( D => n8086, CK => clk, Q => 
                           n6756, QN => n4472);
   registers_reg_13_38_inst : DFF_X1 port map( D => n8085, CK => clk, Q => 
                           n6823, QN => n4473);
   registers_reg_13_37_inst : DFF_X1 port map( D => n8084, CK => clk, Q => 
                           n6890, QN => n4474);
   registers_reg_13_36_inst : DFF_X1 port map( D => n8083, CK => clk, Q => 
                           n6957, QN => n4475);
   registers_reg_13_35_inst : DFF_X1 port map( D => n8082, CK => clk, Q => 
                           n9263, QN => n4476);
   registers_reg_13_34_inst : DFF_X1 port map( D => n8081, CK => clk, Q => 
                           n9331, QN => n4477);
   registers_reg_13_33_inst : DFF_X1 port map( D => n8080, CK => clk, Q => 
                           n9398, QN => n4478);
   registers_reg_13_32_inst : DFF_X1 port map( D => n8079, CK => clk, Q => 
                           n9465, QN => n4479);
   registers_reg_13_31_inst : DFF_X1 port map( D => n8078, CK => clk, Q => 
                           n9533, QN => n4480);
   registers_reg_13_30_inst : DFF_X1 port map( D => n8077, CK => clk, Q => 
                           n9600, QN => n4481);
   registers_reg_13_29_inst : DFF_X1 port map( D => n8076, CK => clk, Q => 
                           n9667, QN => n4482);
   registers_reg_13_28_inst : DFF_X1 port map( D => n8075, CK => clk, Q => 
                           n9734, QN => n4483);
   registers_reg_13_27_inst : DFF_X1 port map( D => n8074, CK => clk, Q => 
                           n9802, QN => n4484);
   registers_reg_13_26_inst : DFF_X1 port map( D => n8073, CK => clk, Q => 
                           n9869, QN => n4485);
   registers_reg_13_25_inst : DFF_X1 port map( D => n8072, CK => clk, Q => 
                           n9936, QN => n4486);
   registers_reg_13_24_inst : DFF_X1 port map( D => n8071, CK => clk, Q => 
                           n10003, QN => n4487);
   registers_reg_13_23_inst : DFF_X1 port map( D => n8070, CK => clk, Q => 
                           n10071, QN => n4488);
   registers_reg_13_22_inst : DFF_X1 port map( D => n8069, CK => clk, Q => 
                           n10138, QN => n4489);
   registers_reg_13_21_inst : DFF_X1 port map( D => n8068, CK => clk, Q => 
                           n10205, QN => n4490);
   registers_reg_13_20_inst : DFF_X1 port map( D => n8067, CK => clk, Q => 
                           n10273, QN => n4491);
   registers_reg_13_19_inst : DFF_X1 port map( D => n8066, CK => clk, Q => 
                           n10340, QN => n4492);
   registers_reg_13_18_inst : DFF_X1 port map( D => n8065, CK => clk, Q => 
                           n10407, QN => n4493);
   registers_reg_13_17_inst : DFF_X1 port map( D => n8064, CK => clk, Q => 
                           n10474, QN => n4494);
   registers_reg_13_16_inst : DFF_X1 port map( D => n8063, CK => clk, Q => 
                           n10542, QN => n4495);
   registers_reg_13_15_inst : DFF_X1 port map( D => n8062, CK => clk, Q => 
                           n10609, QN => n4496);
   registers_reg_13_14_inst : DFF_X1 port map( D => n8061, CK => clk, Q => 
                           n10676, QN => n4497);
   registers_reg_13_13_inst : DFF_X1 port map( D => n8060, CK => clk, Q => 
                           n10743, QN => n4498);
   registers_reg_13_12_inst : DFF_X1 port map( D => n8059, CK => clk, Q => 
                           n10811, QN => n4499);
   registers_reg_13_11_inst : DFF_X1 port map( D => n8058, CK => clk, Q => 
                           n10878, QN => n4500);
   registers_reg_13_10_inst : DFF_X1 port map( D => n8057, CK => clk, Q => 
                           n10945, QN => n4501);
   registers_reg_13_9_inst : DFF_X1 port map( D => n8056, CK => clk, Q => 
                           n11012, QN => n4502);
   registers_reg_13_8_inst : DFF_X1 port map( D => n8055, CK => clk, Q => 
                           n11080, QN => n4503);
   registers_reg_13_7_inst : DFF_X1 port map( D => n8054, CK => clk, Q => 
                           n11147, QN => n4504);
   registers_reg_13_6_inst : DFF_X1 port map( D => n8053, CK => clk, Q => 
                           n11214, QN => n4505);
   registers_reg_13_5_inst : DFF_X1 port map( D => n8052, CK => clk, Q => 
                           n11282, QN => n4506);
   registers_reg_13_4_inst : DFF_X1 port map( D => n8051, CK => clk, Q => 
                           n11349, QN => n4507);
   registers_reg_30_3_inst : DFF_X1 port map( D => n9138, CK => clk, Q => 
                           n18885, QN => n3363);
   registers_reg_30_2_inst : DFF_X1 port map( D => n9137, CK => clk, Q => 
                           n18884, QN => n3364);
   registers_reg_30_1_inst : DFF_X1 port map( D => n9136, CK => clk, Q => 
                           n18883, QN => n3365);
   registers_reg_30_0_inst : DFF_X1 port map( D => n9135, CK => clk, Q => 
                           n18882, QN => n3366);
   registers_reg_12_63_inst : DFF_X1 port map( D => n8046, CK => clk, Q => 
                           n18881, QN => n4517);
   registers_reg_12_62_inst : DFF_X1 port map( D => n8045, CK => clk, Q => 
                           n18880, QN => n4518);
   registers_reg_12_61_inst : DFF_X1 port map( D => n8044, CK => clk, Q => 
                           n18879, QN => n4519);
   registers_reg_12_60_inst : DFF_X1 port map( D => n8043, CK => clk, Q => 
                           n18878, QN => n4520);
   registers_reg_12_59_inst : DFF_X1 port map( D => n8042, CK => clk, Q => 
                           n18877, QN => n4521);
   registers_reg_12_58_inst : DFF_X1 port map( D => n8041, CK => clk, Q => 
                           n18876, QN => n4522);
   registers_reg_12_57_inst : DFF_X1 port map( D => n8040, CK => clk, Q => 
                           n18875, QN => n4523);
   registers_reg_12_56_inst : DFF_X1 port map( D => n8039, CK => clk, Q => 
                           n18874, QN => n4524);
   registers_reg_12_55_inst : DFF_X1 port map( D => n8038, CK => clk, Q => 
                           n18873, QN => n4525);
   registers_reg_12_54_inst : DFF_X1 port map( D => n8037, CK => clk, Q => 
                           n18872, QN => n4526);
   registers_reg_12_53_inst : DFF_X1 port map( D => n8036, CK => clk, Q => 
                           n18871, QN => n4527);
   registers_reg_12_52_inst : DFF_X1 port map( D => n8035, CK => clk, Q => 
                           n18870, QN => n4528);
   registers_reg_12_51_inst : DFF_X1 port map( D => n8034, CK => clk, Q => 
                           n18869, QN => n4529);
   registers_reg_12_50_inst : DFF_X1 port map( D => n8033, CK => clk, Q => 
                           n18868, QN => n4530);
   registers_reg_12_49_inst : DFF_X1 port map( D => n8032, CK => clk, Q => 
                           n18867, QN => n4531);
   registers_reg_12_48_inst : DFF_X1 port map( D => n8031, CK => clk, Q => 
                           n18866, QN => n4532);
   registers_reg_12_47_inst : DFF_X1 port map( D => n8030, CK => clk, Q => 
                           n18865, QN => n4533);
   registers_reg_12_46_inst : DFF_X1 port map( D => n8029, CK => clk, Q => 
                           n18864, QN => n4534);
   registers_reg_12_45_inst : DFF_X1 port map( D => n8028, CK => clk, Q => 
                           n18863, QN => n4535);
   registers_reg_12_44_inst : DFF_X1 port map( D => n8027, CK => clk, Q => 
                           n18862, QN => n4536);
   registers_reg_12_43_inst : DFF_X1 port map( D => n8026, CK => clk, Q => 
                           n18861, QN => n4537);
   registers_reg_12_42_inst : DFF_X1 port map( D => n8025, CK => clk, Q => 
                           n18860, QN => n4538);
   registers_reg_12_41_inst : DFF_X1 port map( D => n8024, CK => clk, Q => 
                           n18859, QN => n4539);
   registers_reg_12_40_inst : DFF_X1 port map( D => n8023, CK => clk, Q => 
                           n18858, QN => n4540);
   registers_reg_12_39_inst : DFF_X1 port map( D => n8022, CK => clk, Q => 
                           n18857, QN => n4541);
   registers_reg_12_38_inst : DFF_X1 port map( D => n8021, CK => clk, Q => 
                           n18856, QN => n4542);
   registers_reg_12_37_inst : DFF_X1 port map( D => n8020, CK => clk, Q => 
                           n18855, QN => n4543);
   registers_reg_12_36_inst : DFF_X1 port map( D => n8019, CK => clk, Q => 
                           n18854, QN => n4544);
   registers_reg_12_35_inst : DFF_X1 port map( D => n8018, CK => clk, Q => 
                           n18853, QN => n4545);
   registers_reg_12_34_inst : DFF_X1 port map( D => n8017, CK => clk, Q => 
                           n18852, QN => n4546);
   registers_reg_12_33_inst : DFF_X1 port map( D => n8016, CK => clk, Q => 
                           n18851, QN => n4547);
   registers_reg_12_32_inst : DFF_X1 port map( D => n8015, CK => clk, Q => 
                           n18850, QN => n4548);
   registers_reg_12_31_inst : DFF_X1 port map( D => n8014, CK => clk, Q => 
                           n18849, QN => n4549);
   registers_reg_12_30_inst : DFF_X1 port map( D => n8013, CK => clk, Q => 
                           n18848, QN => n4550);
   registers_reg_12_29_inst : DFF_X1 port map( D => n8012, CK => clk, Q => 
                           n18847, QN => n4551);
   registers_reg_12_28_inst : DFF_X1 port map( D => n8011, CK => clk, Q => 
                           n18846, QN => n4552);
   registers_reg_12_27_inst : DFF_X1 port map( D => n8010, CK => clk, Q => 
                           n18845, QN => n4553);
   registers_reg_12_26_inst : DFF_X1 port map( D => n8009, CK => clk, Q => 
                           n18844, QN => n4554);
   registers_reg_12_25_inst : DFF_X1 port map( D => n8008, CK => clk, Q => 
                           n18843, QN => n4555);
   registers_reg_12_24_inst : DFF_X1 port map( D => n8007, CK => clk, Q => 
                           n18842, QN => n4556);
   registers_reg_12_23_inst : DFF_X1 port map( D => n8006, CK => clk, Q => 
                           n18841, QN => n4557);
   registers_reg_12_22_inst : DFF_X1 port map( D => n8005, CK => clk, Q => 
                           n18840, QN => n4558);
   registers_reg_12_21_inst : DFF_X1 port map( D => n8004, CK => clk, Q => 
                           n18839, QN => n4559);
   registers_reg_12_20_inst : DFF_X1 port map( D => n8003, CK => clk, Q => 
                           n18838, QN => n4560);
   registers_reg_12_19_inst : DFF_X1 port map( D => n8002, CK => clk, Q => 
                           n18837, QN => n4561);
   registers_reg_12_18_inst : DFF_X1 port map( D => n8001, CK => clk, Q => 
                           n18836, QN => n4562);
   registers_reg_12_17_inst : DFF_X1 port map( D => n8000, CK => clk, Q => 
                           n18835, QN => n4563);
   registers_reg_12_16_inst : DFF_X1 port map( D => n7999, CK => clk, Q => 
                           n18834, QN => n4564);
   registers_reg_12_15_inst : DFF_X1 port map( D => n7998, CK => clk, Q => 
                           n18833, QN => n4565);
   registers_reg_12_14_inst : DFF_X1 port map( D => n7997, CK => clk, Q => 
                           n18832, QN => n4566);
   registers_reg_12_13_inst : DFF_X1 port map( D => n7996, CK => clk, Q => 
                           n18831, QN => n4567);
   registers_reg_12_12_inst : DFF_X1 port map( D => n7995, CK => clk, Q => 
                           n18830, QN => n4568);
   registers_reg_12_11_inst : DFF_X1 port map( D => n7994, CK => clk, Q => 
                           n18829, QN => n4569);
   registers_reg_12_10_inst : DFF_X1 port map( D => n7993, CK => clk, Q => 
                           n18828, QN => n4570);
   registers_reg_12_9_inst : DFF_X1 port map( D => n7992, CK => clk, Q => 
                           n18827, QN => n4571);
   registers_reg_12_8_inst : DFF_X1 port map( D => n7991, CK => clk, Q => 
                           n18826, QN => n4572);
   registers_reg_12_7_inst : DFF_X1 port map( D => n7990, CK => clk, Q => 
                           n18825, QN => n4573);
   registers_reg_12_6_inst : DFF_X1 port map( D => n7989, CK => clk, Q => 
                           n18824, QN => n4574);
   registers_reg_12_5_inst : DFF_X1 port map( D => n7988, CK => clk, Q => 
                           n18823, QN => n4575);
   registers_reg_12_4_inst : DFF_X1 port map( D => n7987, CK => clk, Q => 
                           n18822, QN => n4576);
   registers_reg_6_3_inst : DFF_X1 port map( D => n7602, CK => clk, Q => n11366
                           , QN => n4984);
   registers_reg_6_2_inst : DFF_X1 port map( D => n7601, CK => clk, Q => n11433
                           , QN => n4985);
   registers_reg_6_1_inst : DFF_X1 port map( D => n7600, CK => clk, Q => n11501
                           , QN => n4986);
   registers_reg_6_0_inst : DFF_X1 port map( D => n7599, CK => clk, Q => n11593
                           , QN => n4987);
   registers_reg_5_3_inst : DFF_X1 port map( D => n7538, CK => clk, Q => n11363
                           , QN => n5050);
   registers_reg_5_2_inst : DFF_X1 port map( D => n7537, CK => clk, Q => n11430
                           , QN => n5051);
   registers_reg_5_1_inst : DFF_X1 port map( D => n7536, CK => clk, Q => n11498
                           , QN => n5052);
   registers_reg_5_0_inst : DFF_X1 port map( D => n7535, CK => clk, Q => n11585
                           , QN => n5053);
   registers_reg_7_3_inst : DFF_X1 port map( D => n7666, CK => clk, Q => n11419
                           , QN => n4918);
   registers_reg_7_2_inst : DFF_X1 port map( D => n7665, CK => clk, Q => n11486
                           , QN => n4919);
   registers_reg_7_1_inst : DFF_X1 port map( D => n7664, CK => clk, Q => n11554
                           , QN => n4920);
   registers_reg_7_0_inst : DFF_X1 port map( D => n7663, CK => clk, Q => n11719
                           , QN => n4921);
   registers_reg_25_3_inst : DFF_X1 port map( D => n8818, CK => clk, Q => 
                           n11371, QN => n3701);
   registers_reg_25_2_inst : DFF_X1 port map( D => n8817, CK => clk, Q => 
                           n11439, QN => n3702);
   registers_reg_25_1_inst : DFF_X1 port map( D => n8816, CK => clk, Q => 
                           n11506, QN => n3703);
   registers_reg_25_0_inst : DFF_X1 port map( D => n8815, CK => clk, Q => 
                           n11605, QN => n3704);
   registers_reg_17_3_inst : DFF_X1 port map( D => n8306, CK => clk, Q => 
                           n18821, QN => n4239);
   registers_reg_17_2_inst : DFF_X1 port map( D => n8305, CK => clk, Q => 
                           n18820, QN => n4240);
   registers_reg_17_1_inst : DFF_X1 port map( D => n8304, CK => clk, Q => 
                           n18819, QN => n4241);
   registers_reg_17_0_inst : DFF_X1 port map( D => n8303, CK => clk, Q => 
                           n18818, QN => n4242);
   registers_reg_20_3_inst : DFF_X1 port map( D => n8498, CK => clk, Q => 
                           n11372, QN => n4034);
   registers_reg_20_2_inst : DFF_X1 port map( D => n8497, CK => clk, Q => 
                           n11440, QN => n4035);
   registers_reg_20_1_inst : DFF_X1 port map( D => n8496, CK => clk, Q => 
                           n11507, QN => n4036);
   registers_reg_20_0_inst : DFF_X1 port map( D => n8495, CK => clk, Q => 
                           n11606, QN => n4037);
   registers_reg_31_3_inst : DFF_X1 port map( D => n9202, CK => clk, Q => 
                           n11369, QN => n3289);
   registers_reg_31_2_inst : DFF_X1 port map( D => n9201, CK => clk, Q => 
                           n11437, QN => n3291);
   registers_reg_31_1_inst : DFF_X1 port map( D => n9200, CK => clk, Q => 
                           n11504, QN => n3293);
   registers_reg_31_0_inst : DFF_X1 port map( D => n9199, CK => clk, Q => 
                           n11599, QN => n3295);
   registers_reg_27_3_inst : DFF_X1 port map( D => n8946, CK => clk, Q => 
                           n11415, QN => n3566);
   registers_reg_27_2_inst : DFF_X1 port map( D => n8945, CK => clk, Q => 
                           n11482, QN => n3567);
   registers_reg_27_1_inst : DFF_X1 port map( D => n8944, CK => clk, Q => 
                           n11550, QN => n3568);
   registers_reg_27_0_inst : DFF_X1 port map( D => n8943, CK => clk, Q => 
                           n11704, QN => n3569);
   registers_reg_19_3_inst : DFF_X1 port map( D => n8434, CK => clk, Q => 
                           n11364, QN => n4100);
   registers_reg_19_2_inst : DFF_X1 port map( D => n8433, CK => clk, Q => 
                           n11431, QN => n4101);
   registers_reg_19_1_inst : DFF_X1 port map( D => n8432, CK => clk, Q => 
                           n11499, QN => n4102);
   registers_reg_19_0_inst : DFF_X1 port map( D => n8431, CK => clk, Q => 
                           n11586, QN => n4103);
   registers_reg_29_3_inst : DFF_X1 port map( D => n9074, CK => clk, Q => 
                           n18817, QN => n3431);
   registers_reg_29_2_inst : DFF_X1 port map( D => n9073, CK => clk, Q => 
                           n18816, QN => n3432);
   registers_reg_29_1_inst : DFF_X1 port map( D => n9072, CK => clk, Q => 
                           n18815, QN => n3433);
   registers_reg_29_0_inst : DFF_X1 port map( D => n9071, CK => clk, Q => 
                           n18814, QN => n3434);
   registers_reg_1_63_inst : DFF_X1 port map( D => n7342, CK => clk, Q => 
                           n18813, QN => n5257);
   registers_reg_1_62_inst : DFF_X1 port map( D => n7341, CK => clk, Q => 
                           n18812, QN => n5258);
   registers_reg_1_61_inst : DFF_X1 port map( D => n7340, CK => clk, Q => 
                           n18811, QN => n5259);
   registers_reg_1_60_inst : DFF_X1 port map( D => n7339, CK => clk, Q => 
                           n18810, QN => n5260);
   registers_reg_1_59_inst : DFF_X1 port map( D => n7338, CK => clk, Q => 
                           n18809, QN => n5261);
   registers_reg_1_58_inst : DFF_X1 port map( D => n7337, CK => clk, Q => 
                           n18808, QN => n5262);
   registers_reg_1_57_inst : DFF_X1 port map( D => n7336, CK => clk, Q => 
                           n18807, QN => n5263);
   registers_reg_1_56_inst : DFF_X1 port map( D => n7335, CK => clk, Q => 
                           n18806, QN => n5264);
   registers_reg_1_55_inst : DFF_X1 port map( D => n7334, CK => clk, Q => 
                           n18805, QN => n5265);
   registers_reg_1_54_inst : DFF_X1 port map( D => n7333, CK => clk, Q => 
                           n18804, QN => n5266);
   registers_reg_1_53_inst : DFF_X1 port map( D => n7332, CK => clk, Q => 
                           n18803, QN => n5267);
   registers_reg_1_52_inst : DFF_X1 port map( D => n7331, CK => clk, Q => 
                           n18802, QN => n5268);
   registers_reg_1_51_inst : DFF_X1 port map( D => n7330, CK => clk, Q => 
                           n18801, QN => n5269);
   registers_reg_1_50_inst : DFF_X1 port map( D => n7329, CK => clk, Q => 
                           n18800, QN => n5270);
   registers_reg_1_49_inst : DFF_X1 port map( D => n7328, CK => clk, Q => 
                           n18799, QN => n5271);
   registers_reg_1_48_inst : DFF_X1 port map( D => n7327, CK => clk, Q => 
                           n18798, QN => n5272);
   registers_reg_1_47_inst : DFF_X1 port map( D => n7326, CK => clk, Q => 
                           n18797, QN => n5273);
   registers_reg_1_46_inst : DFF_X1 port map( D => n7325, CK => clk, Q => 
                           n18796, QN => n5274);
   registers_reg_1_45_inst : DFF_X1 port map( D => n7324, CK => clk, Q => 
                           n18795, QN => n5275);
   registers_reg_1_44_inst : DFF_X1 port map( D => n7323, CK => clk, Q => 
                           n18794, QN => n5276);
   registers_reg_1_43_inst : DFF_X1 port map( D => n7322, CK => clk, Q => 
                           n18793, QN => n5277);
   registers_reg_1_42_inst : DFF_X1 port map( D => n7321, CK => clk, Q => 
                           n18792, QN => n5278);
   registers_reg_1_41_inst : DFF_X1 port map( D => n7320, CK => clk, Q => 
                           n18791, QN => n5279);
   registers_reg_1_40_inst : DFF_X1 port map( D => n7319, CK => clk, Q => 
                           n18790, QN => n5280);
   registers_reg_1_39_inst : DFF_X1 port map( D => n7318, CK => clk, Q => 
                           n18789, QN => n5281);
   registers_reg_1_38_inst : DFF_X1 port map( D => n7317, CK => clk, Q => 
                           n18788, QN => n5282);
   registers_reg_1_37_inst : DFF_X1 port map( D => n7316, CK => clk, Q => 
                           n18787, QN => n5283);
   registers_reg_1_36_inst : DFF_X1 port map( D => n7315, CK => clk, Q => 
                           n18786, QN => n5284);
   registers_reg_1_35_inst : DFF_X1 port map( D => n7314, CK => clk, Q => 
                           n18785, QN => n5285);
   registers_reg_1_34_inst : DFF_X1 port map( D => n7313, CK => clk, Q => 
                           n18784, QN => n5286);
   registers_reg_1_33_inst : DFF_X1 port map( D => n7312, CK => clk, Q => 
                           n18783, QN => n5287);
   registers_reg_1_32_inst : DFF_X1 port map( D => n7311, CK => clk, Q => 
                           n18782, QN => n5288);
   registers_reg_1_31_inst : DFF_X1 port map( D => n7310, CK => clk, Q => 
                           n18781, QN => n5289);
   registers_reg_1_30_inst : DFF_X1 port map( D => n7309, CK => clk, Q => 
                           n18780, QN => n5290);
   registers_reg_1_29_inst : DFF_X1 port map( D => n7308, CK => clk, Q => 
                           n18779, QN => n5291);
   registers_reg_1_28_inst : DFF_X1 port map( D => n7307, CK => clk, Q => 
                           n18778, QN => n5355);
   registers_reg_1_27_inst : DFF_X1 port map( D => n7306, CK => clk, Q => 
                           n18777, QN => n5356);
   registers_reg_1_26_inst : DFF_X1 port map( D => n7305, CK => clk, Q => 
                           n18776, QN => n5357);
   registers_reg_1_25_inst : DFF_X1 port map( D => n7304, CK => clk, Q => 
                           n18775, QN => n5359);
   registers_reg_1_24_inst : DFF_X1 port map( D => n7303, CK => clk, Q => 
                           n18774, QN => n5424);
   registers_reg_1_23_inst : DFF_X1 port map( D => n7302, CK => clk, Q => 
                           n18773, QN => n5426);
   registers_reg_1_22_inst : DFF_X1 port map( D => n7301, CK => clk, Q => 
                           n18772, QN => n5491);
   registers_reg_1_21_inst : DFF_X1 port map( D => n7300, CK => clk, Q => 
                           n18771, QN => n5492);
   registers_reg_1_20_inst : DFF_X1 port map( D => n7299, CK => clk, Q => 
                           n18770, QN => n5494);
   registers_reg_1_19_inst : DFF_X1 port map( D => n7298, CK => clk, Q => 
                           n18769, QN => n5559);
   registers_reg_1_18_inst : DFF_X1 port map( D => n7297, CK => clk, Q => 
                           n18768, QN => n5560);
   registers_reg_1_17_inst : DFF_X1 port map( D => n7296, CK => clk, Q => 
                           n18767, QN => n5562);
   registers_reg_1_16_inst : DFF_X1 port map( D => n7295, CK => clk, Q => 
                           n18766, QN => n5627);
   registers_reg_1_15_inst : DFF_X1 port map( D => n7294, CK => clk, Q => 
                           n18765, QN => n5629);
   registers_reg_1_14_inst : DFF_X1 port map( D => n7293, CK => clk, Q => 
                           n18764, QN => n5694);
   registers_reg_1_13_inst : DFF_X1 port map( D => n7292, CK => clk, Q => 
                           n18763, QN => n5695);
   registers_reg_1_12_inst : DFF_X1 port map( D => n7291, CK => clk, Q => 
                           n18762, QN => n5696);
   registers_reg_1_11_inst : DFF_X1 port map( D => n7290, CK => clk, Q => 
                           n18761, QN => n5698);
   registers_reg_1_10_inst : DFF_X1 port map( D => n7289, CK => clk, Q => 
                           n18760, QN => n5763);
   registers_reg_1_9_inst : DFF_X1 port map( D => n7288, CK => clk, Q => n18759
                           , QN => n5764);
   registers_reg_1_8_inst : DFF_X1 port map( D => n7287, CK => clk, Q => n18758
                           , QN => n5765);
   registers_reg_1_7_inst : DFF_X1 port map( D => n7286, CK => clk, Q => n18757
                           , QN => n5766);
   registers_reg_1_6_inst : DFF_X1 port map( D => n7285, CK => clk, Q => n18756
                           , QN => n5767);
   registers_reg_1_5_inst : DFF_X1 port map( D => n7284, CK => clk, Q => n18755
                           , QN => n5769);
   registers_reg_1_4_inst : DFF_X1 port map( D => n7283, CK => clk, Q => n18754
                           , QN => n5835);
   registers_reg_16_63_inst : DFF_X1 port map( D => n8302, CK => clk, Q => 
                           n3018, QN => n4246);
   registers_reg_16_62_inst : DFF_X1 port map( D => n8301, CK => clk, Q => 
                           n3258, QN => n4247);
   registers_reg_16_61_inst : DFF_X1 port map( D => n8300, CK => clk, Q => 
                           n4175, QN => n4248);
   registers_reg_16_60_inst : DFF_X1 port map( D => n8299, CK => clk, Q => 
                           n5300, QN => n4249);
   registers_reg_16_59_inst : DFF_X1 port map( D => n8298, CK => clk, Q => 
                           n5370, QN => n4250);
   registers_reg_16_58_inst : DFF_X1 port map( D => n8297, CK => clk, Q => 
                           n5438, QN => n4251);
   registers_reg_16_57_inst : DFF_X1 port map( D => n8296, CK => clk, Q => 
                           n5507, QN => n4252);
   registers_reg_16_56_inst : DFF_X1 port map( D => n8295, CK => clk, Q => 
                           n5576, QN => n4253);
   registers_reg_16_55_inst : DFF_X1 port map( D => n8294, CK => clk, Q => 
                           n5644, QN => n4254);
   registers_reg_16_54_inst : DFF_X1 port map( D => n8293, CK => clk, Q => 
                           n5714, QN => n4255);
   registers_reg_16_53_inst : DFF_X1 port map( D => n8292, CK => clk, Q => 
                           n5786, QN => n4256);
   registers_reg_16_52_inst : DFF_X1 port map( D => n8291, CK => clk, Q => 
                           n5853, QN => n4257);
   registers_reg_16_51_inst : DFF_X1 port map( D => n8290, CK => clk, Q => 
                           n5920, QN => n4258);
   registers_reg_16_50_inst : DFF_X1 port map( D => n8289, CK => clk, Q => 
                           n5988, QN => n4259);
   registers_reg_16_49_inst : DFF_X1 port map( D => n8288, CK => clk, Q => 
                           n6056, QN => n4260);
   registers_reg_16_48_inst : DFF_X1 port map( D => n8287, CK => clk, Q => 
                           n6122, QN => n4261);
   registers_reg_16_47_inst : DFF_X1 port map( D => n8286, CK => clk, Q => 
                           n6188, QN => n4262);
   registers_reg_16_46_inst : DFF_X1 port map( D => n8285, CK => clk, Q => 
                           n6254, QN => n4263);
   registers_reg_16_45_inst : DFF_X1 port map( D => n8284, CK => clk, Q => 
                           n6320, QN => n4264);
   registers_reg_16_44_inst : DFF_X1 port map( D => n8283, CK => clk, Q => 
                           n6386, QN => n4265);
   registers_reg_16_43_inst : DFF_X1 port map( D => n8282, CK => clk, Q => 
                           n6452, QN => n4266);
   registers_reg_16_42_inst : DFF_X1 port map( D => n8281, CK => clk, Q => 
                           n6518, QN => n4267);
   registers_reg_16_41_inst : DFF_X1 port map( D => n8280, CK => clk, Q => 
                           n6584, QN => n4268);
   registers_reg_16_40_inst : DFF_X1 port map( D => n8279, CK => clk, Q => 
                           n6651, QN => n4269);
   registers_reg_16_39_inst : DFF_X1 port map( D => n8278, CK => clk, Q => 
                           n6718, QN => n4270);
   registers_reg_16_38_inst : DFF_X1 port map( D => n8277, CK => clk, Q => 
                           n6785, QN => n4271);
   registers_reg_16_37_inst : DFF_X1 port map( D => n8276, CK => clk, Q => 
                           n6852, QN => n4272);
   registers_reg_16_36_inst : DFF_X1 port map( D => n8275, CK => clk, Q => 
                           n6919, QN => n4273);
   registers_reg_16_35_inst : DFF_X1 port map( D => n8274, CK => clk, Q => 
                           n6986, QN => n4274);
   registers_reg_16_34_inst : DFF_X1 port map( D => n8273, CK => clk, Q => 
                           n9293, QN => n4275);
   registers_reg_16_33_inst : DFF_X1 port map( D => n8272, CK => clk, Q => 
                           n9360, QN => n4276);
   registers_reg_16_32_inst : DFF_X1 port map( D => n8271, CK => clk, Q => 
                           n9428, QN => n4277);
   registers_reg_16_31_inst : DFF_X1 port map( D => n8270, CK => clk, Q => 
                           n9495, QN => n4278);
   registers_reg_16_30_inst : DFF_X1 port map( D => n8269, CK => clk, Q => 
                           n9562, QN => n4279);
   registers_reg_16_29_inst : DFF_X1 port map( D => n8268, CK => clk, Q => 
                           n9629, QN => n4280);
   registers_reg_16_28_inst : DFF_X1 port map( D => n8267, CK => clk, Q => 
                           n9697, QN => n4281);
   registers_reg_16_27_inst : DFF_X1 port map( D => n8266, CK => clk, Q => 
                           n9764, QN => n4282);
   registers_reg_16_26_inst : DFF_X1 port map( D => n8265, CK => clk, Q => 
                           n9831, QN => n4283);
   registers_reg_16_25_inst : DFF_X1 port map( D => n8264, CK => clk, Q => 
                           n9898, QN => n4284);
   registers_reg_16_24_inst : DFF_X1 port map( D => n8263, CK => clk, Q => 
                           n9966, QN => n4285);
   registers_reg_16_23_inst : DFF_X1 port map( D => n8262, CK => clk, Q => 
                           n10033, QN => n4286);
   registers_reg_16_22_inst : DFF_X1 port map( D => n8261, CK => clk, Q => 
                           n10100, QN => n4287);
   registers_reg_16_21_inst : DFF_X1 port map( D => n8260, CK => clk, Q => 
                           n10168, QN => n4288);
   registers_reg_16_20_inst : DFF_X1 port map( D => n8259, CK => clk, Q => 
                           n10235, QN => n4289);
   registers_reg_16_19_inst : DFF_X1 port map( D => n8258, CK => clk, Q => 
                           n10302, QN => n4290);
   registers_reg_16_18_inst : DFF_X1 port map( D => n8257, CK => clk, Q => 
                           n10369, QN => n4291);
   registers_reg_16_17_inst : DFF_X1 port map( D => n8256, CK => clk, Q => 
                           n10437, QN => n4292);
   registers_reg_16_16_inst : DFF_X1 port map( D => n8255, CK => clk, Q => 
                           n10504, QN => n4293);
   registers_reg_16_15_inst : DFF_X1 port map( D => n8254, CK => clk, Q => 
                           n10571, QN => n4294);
   registers_reg_16_14_inst : DFF_X1 port map( D => n8253, CK => clk, Q => 
                           n10638, QN => n4295);
   registers_reg_16_13_inst : DFF_X1 port map( D => n8252, CK => clk, Q => 
                           n10706, QN => n4296);
   registers_reg_16_12_inst : DFF_X1 port map( D => n8251, CK => clk, Q => 
                           n10773, QN => n4297);
   registers_reg_16_11_inst : DFF_X1 port map( D => n8250, CK => clk, Q => 
                           n10840, QN => n4298);
   registers_reg_16_10_inst : DFF_X1 port map( D => n8249, CK => clk, Q => 
                           n10908, QN => n4299);
   registers_reg_16_9_inst : DFF_X1 port map( D => n8248, CK => clk, Q => 
                           n10975, QN => n4300);
   registers_reg_16_8_inst : DFF_X1 port map( D => n8247, CK => clk, Q => 
                           n11042, QN => n4301);
   registers_reg_16_7_inst : DFF_X1 port map( D => n8246, CK => clk, Q => 
                           n11109, QN => n4302);
   registers_reg_16_6_inst : DFF_X1 port map( D => n8245, CK => clk, Q => 
                           n11177, QN => n4303);
   registers_reg_16_5_inst : DFF_X1 port map( D => n8244, CK => clk, Q => 
                           n11244, QN => n4304);
   registers_reg_16_4_inst : DFF_X1 port map( D => n8243, CK => clk, Q => 
                           n11311, QN => n4305);
   registers_reg_23_3_inst : DFF_X1 port map( D => n8690, CK => clk, Q => 
                           n18753, QN => n3833);
   registers_reg_23_2_inst : DFF_X1 port map( D => n8689, CK => clk, Q => 
                           n18752, QN => n3834);
   registers_reg_23_1_inst : DFF_X1 port map( D => n8688, CK => clk, Q => 
                           n18751, QN => n3835);
   registers_reg_23_0_inst : DFF_X1 port map( D => n8687, CK => clk, Q => 
                           n18750, QN => n3836);
   registers_reg_28_63_inst : DFF_X1 port map( D => n9070, CK => clk, Q => 
                           n18749, QN => n3439);
   registers_reg_28_62_inst : DFF_X1 port map( D => n9069, CK => clk, Q => 
                           n18748, QN => n3440);
   registers_reg_28_61_inst : DFF_X1 port map( D => n9068, CK => clk, Q => 
                           n18747, QN => n3441);
   registers_reg_28_60_inst : DFF_X1 port map( D => n9067, CK => clk, Q => 
                           n18746, QN => n3442);
   registers_reg_28_59_inst : DFF_X1 port map( D => n9066, CK => clk, Q => 
                           n18745, QN => n3443);
   registers_reg_28_58_inst : DFF_X1 port map( D => n9065, CK => clk, Q => 
                           n18744, QN => n3444);
   registers_reg_28_57_inst : DFF_X1 port map( D => n9064, CK => clk, Q => 
                           n18743, QN => n3445);
   registers_reg_28_56_inst : DFF_X1 port map( D => n9063, CK => clk, Q => 
                           n18742, QN => n3446);
   registers_reg_28_55_inst : DFF_X1 port map( D => n9062, CK => clk, Q => 
                           n18741, QN => n3447);
   registers_reg_28_54_inst : DFF_X1 port map( D => n9061, CK => clk, Q => 
                           n18740, QN => n3448);
   registers_reg_28_53_inst : DFF_X1 port map( D => n9060, CK => clk, Q => 
                           n18739, QN => n3449);
   registers_reg_28_52_inst : DFF_X1 port map( D => n9059, CK => clk, Q => 
                           n18738, QN => n3450);
   registers_reg_28_51_inst : DFF_X1 port map( D => n9058, CK => clk, Q => 
                           n18737, QN => n3451);
   registers_reg_28_50_inst : DFF_X1 port map( D => n9057, CK => clk, Q => 
                           n18736, QN => n3452);
   registers_reg_28_49_inst : DFF_X1 port map( D => n9056, CK => clk, Q => 
                           n18735, QN => n3453);
   registers_reg_28_48_inst : DFF_X1 port map( D => n9055, CK => clk, Q => 
                           n18734, QN => n3454);
   registers_reg_28_47_inst : DFF_X1 port map( D => n9054, CK => clk, Q => 
                           n18733, QN => n3455);
   registers_reg_28_46_inst : DFF_X1 port map( D => n9053, CK => clk, Q => 
                           n18732, QN => n3456);
   registers_reg_28_45_inst : DFF_X1 port map( D => n9052, CK => clk, Q => 
                           n18731, QN => n3457);
   registers_reg_28_44_inst : DFF_X1 port map( D => n9051, CK => clk, Q => 
                           n18730, QN => n3458);
   registers_reg_28_43_inst : DFF_X1 port map( D => n9050, CK => clk, Q => 
                           n18729, QN => n3459);
   registers_reg_28_42_inst : DFF_X1 port map( D => n9049, CK => clk, Q => 
                           n18728, QN => n3460);
   registers_reg_28_41_inst : DFF_X1 port map( D => n9048, CK => clk, Q => 
                           n18727, QN => n3461);
   registers_reg_28_40_inst : DFF_X1 port map( D => n9047, CK => clk, Q => 
                           n18726, QN => n3462);
   registers_reg_28_39_inst : DFF_X1 port map( D => n9046, CK => clk, Q => 
                           n18725, QN => n3463);
   registers_reg_28_38_inst : DFF_X1 port map( D => n9045, CK => clk, Q => 
                           n18724, QN => n3464);
   registers_reg_28_37_inst : DFF_X1 port map( D => n9044, CK => clk, Q => 
                           n18723, QN => n3465);
   registers_reg_28_36_inst : DFF_X1 port map( D => n9043, CK => clk, Q => 
                           n18722, QN => n3466);
   registers_reg_28_35_inst : DFF_X1 port map( D => n9042, CK => clk, Q => 
                           n18721, QN => n3467);
   registers_reg_28_34_inst : DFF_X1 port map( D => n9041, CK => clk, Q => 
                           n18720, QN => n3468);
   registers_reg_28_33_inst : DFF_X1 port map( D => n9040, CK => clk, Q => 
                           n18719, QN => n3469);
   registers_reg_28_32_inst : DFF_X1 port map( D => n9039, CK => clk, Q => 
                           n18718, QN => n3470);
   registers_reg_28_31_inst : DFF_X1 port map( D => n9038, CK => clk, Q => 
                           n18717, QN => n3471);
   registers_reg_28_30_inst : DFF_X1 port map( D => n9037, CK => clk, Q => 
                           n18716, QN => n3472);
   registers_reg_28_29_inst : DFF_X1 port map( D => n9036, CK => clk, Q => 
                           n18715, QN => n3473);
   registers_reg_28_28_inst : DFF_X1 port map( D => n9035, CK => clk, Q => 
                           n18714, QN => n3474);
   registers_reg_28_27_inst : DFF_X1 port map( D => n9034, CK => clk, Q => 
                           n18713, QN => n3475);
   registers_reg_28_26_inst : DFF_X1 port map( D => n9033, CK => clk, Q => 
                           n18712, QN => n3476);
   registers_reg_28_25_inst : DFF_X1 port map( D => n9032, CK => clk, Q => 
                           n18711, QN => n3477);
   registers_reg_28_24_inst : DFF_X1 port map( D => n9031, CK => clk, Q => 
                           n18710, QN => n3478);
   registers_reg_28_23_inst : DFF_X1 port map( D => n9030, CK => clk, Q => 
                           n18709, QN => n3479);
   registers_reg_28_22_inst : DFF_X1 port map( D => n9029, CK => clk, Q => 
                           n18708, QN => n3480);
   registers_reg_28_21_inst : DFF_X1 port map( D => n9028, CK => clk, Q => 
                           n18707, QN => n3481);
   registers_reg_28_20_inst : DFF_X1 port map( D => n9027, CK => clk, Q => 
                           n18706, QN => n3482);
   registers_reg_28_19_inst : DFF_X1 port map( D => n9026, CK => clk, Q => 
                           n18705, QN => n3483);
   registers_reg_28_18_inst : DFF_X1 port map( D => n9025, CK => clk, Q => 
                           n18704, QN => n3484);
   registers_reg_28_17_inst : DFF_X1 port map( D => n9024, CK => clk, Q => 
                           n18703, QN => n3485);
   registers_reg_28_16_inst : DFF_X1 port map( D => n9023, CK => clk, Q => 
                           n18702, QN => n3486);
   registers_reg_28_15_inst : DFF_X1 port map( D => n9022, CK => clk, Q => 
                           n18701, QN => n3487);
   registers_reg_28_14_inst : DFF_X1 port map( D => n9021, CK => clk, Q => 
                           n18700, QN => n3488);
   registers_reg_28_13_inst : DFF_X1 port map( D => n9020, CK => clk, Q => 
                           n18699, QN => n3489);
   registers_reg_28_12_inst : DFF_X1 port map( D => n9019, CK => clk, Q => 
                           n18698, QN => n3490);
   registers_reg_28_11_inst : DFF_X1 port map( D => n9018, CK => clk, Q => 
                           n18697, QN => n3491);
   registers_reg_28_10_inst : DFF_X1 port map( D => n9017, CK => clk, Q => 
                           n18696, QN => n3492);
   registers_reg_28_9_inst : DFF_X1 port map( D => n9016, CK => clk, Q => 
                           n18695, QN => n3493);
   registers_reg_28_8_inst : DFF_X1 port map( D => n9015, CK => clk, Q => 
                           n18694, QN => n3494);
   registers_reg_28_7_inst : DFF_X1 port map( D => n9014, CK => clk, Q => 
                           n18693, QN => n3495);
   registers_reg_28_6_inst : DFF_X1 port map( D => n9013, CK => clk, Q => 
                           n18692, QN => n3496);
   registers_reg_28_5_inst : DFF_X1 port map( D => n9012, CK => clk, Q => 
                           n18691, QN => n3497);
   registers_reg_28_4_inst : DFF_X1 port map( D => n9011, CK => clk, Q => 
                           n18690, QN => n3498);
   registers_reg_10_63_inst : DFF_X1 port map( D => n7918, CK => clk, Q => 
                           n3164, QN => n4654);
   registers_reg_10_62_inst : DFF_X1 port map( D => n7917, CK => clk, Q => 
                           n3437, QN => n4655);
   registers_reg_10_61_inst : DFF_X1 port map( D => n7916, CK => clk, Q => 
                           n4719, QN => n4656);
   registers_reg_10_60_inst : DFF_X1 port map( D => n7915, CK => clk, Q => 
                           n5332, QN => n4657);
   registers_reg_10_59_inst : DFF_X1 port map( D => n7914, CK => clk, Q => 
                           n5402, QN => n4658);
   registers_reg_10_58_inst : DFF_X1 port map( D => n7913, CK => clk, Q => 
                           n5470, QN => n4659);
   registers_reg_10_57_inst : DFF_X1 port map( D => n7912, CK => clk, Q => 
                           n5539, QN => n4660);
   registers_reg_10_56_inst : DFF_X1 port map( D => n7911, CK => clk, Q => 
                           n5608, QN => n4661);
   registers_reg_10_55_inst : DFF_X1 port map( D => n7910, CK => clk, Q => 
                           n5676, QN => n4662);
   registers_reg_10_54_inst : DFF_X1 port map( D => n7909, CK => clk, Q => 
                           n5746, QN => n4663);
   registers_reg_10_53_inst : DFF_X1 port map( D => n7908, CK => clk, Q => 
                           n5818, QN => n4664);
   registers_reg_10_52_inst : DFF_X1 port map( D => n7907, CK => clk, Q => 
                           n5885, QN => n4665);
   registers_reg_10_51_inst : DFF_X1 port map( D => n7906, CK => clk, Q => 
                           n5952, QN => n4666);
   registers_reg_10_50_inst : DFF_X1 port map( D => n7905, CK => clk, Q => 
                           n6020, QN => n4667);
   registers_reg_10_49_inst : DFF_X1 port map( D => n7904, CK => clk, Q => 
                           n6088, QN => n4668);
   registers_reg_10_48_inst : DFF_X1 port map( D => n7903, CK => clk, Q => 
                           n6154, QN => n4669);
   registers_reg_10_47_inst : DFF_X1 port map( D => n7902, CK => clk, Q => 
                           n6220, QN => n4670);
   registers_reg_10_46_inst : DFF_X1 port map( D => n7901, CK => clk, Q => 
                           n6286, QN => n4671);
   registers_reg_10_45_inst : DFF_X1 port map( D => n7900, CK => clk, Q => 
                           n6352, QN => n4672);
   registers_reg_10_44_inst : DFF_X1 port map( D => n7899, CK => clk, Q => 
                           n6418, QN => n4673);
   registers_reg_10_43_inst : DFF_X1 port map( D => n7898, CK => clk, Q => 
                           n6484, QN => n4674);
   registers_reg_10_42_inst : DFF_X1 port map( D => n7897, CK => clk, Q => 
                           n6550, QN => n4675);
   registers_reg_10_41_inst : DFF_X1 port map( D => n7896, CK => clk, Q => 
                           n6616, QN => n4676);
   registers_reg_10_40_inst : DFF_X1 port map( D => n7895, CK => clk, Q => 
                           n6683, QN => n4677);
   registers_reg_10_39_inst : DFF_X1 port map( D => n7894, CK => clk, Q => 
                           n6751, QN => n4678);
   registers_reg_10_38_inst : DFF_X1 port map( D => n7893, CK => clk, Q => 
                           n6818, QN => n4679);
   registers_reg_10_37_inst : DFF_X1 port map( D => n7892, CK => clk, Q => 
                           n6885, QN => n4680);
   registers_reg_10_36_inst : DFF_X1 port map( D => n7891, CK => clk, Q => 
                           n6952, QN => n4681);
   registers_reg_10_35_inst : DFF_X1 port map( D => n7890, CK => clk, Q => 
                           n7018, QN => n4682);
   registers_reg_10_34_inst : DFF_X1 port map( D => n7889, CK => clk, Q => 
                           n9326, QN => n4683);
   registers_reg_10_33_inst : DFF_X1 port map( D => n7888, CK => clk, Q => 
                           n9393, QN => n4684);
   registers_reg_10_32_inst : DFF_X1 port map( D => n7887, CK => clk, Q => 
                           n9460, QN => n4685);
   registers_reg_10_31_inst : DFF_X1 port map( D => n7886, CK => clk, Q => 
                           n9527, QN => n4686);
   registers_reg_10_30_inst : DFF_X1 port map( D => n7885, CK => clk, Q => 
                           n9595, QN => n4687);
   registers_reg_10_29_inst : DFF_X1 port map( D => n7884, CK => clk, Q => 
                           n9662, QN => n4688);
   registers_reg_10_28_inst : DFF_X1 port map( D => n7883, CK => clk, Q => 
                           n9729, QN => n4689);
   registers_reg_10_27_inst : DFF_X1 port map( D => n7882, CK => clk, Q => 
                           n9797, QN => n4690);
   registers_reg_10_26_inst : DFF_X1 port map( D => n7881, CK => clk, Q => 
                           n9864, QN => n4691);
   registers_reg_10_25_inst : DFF_X1 port map( D => n7880, CK => clk, Q => 
                           n9931, QN => n4692);
   registers_reg_10_24_inst : DFF_X1 port map( D => n7879, CK => clk, Q => 
                           n9998, QN => n4693);
   registers_reg_10_23_inst : DFF_X1 port map( D => n7878, CK => clk, Q => 
                           n10066, QN => n4694);
   registers_reg_10_22_inst : DFF_X1 port map( D => n7877, CK => clk, Q => 
                           n10133, QN => n4695);
   registers_reg_10_21_inst : DFF_X1 port map( D => n7876, CK => clk, Q => 
                           n10200, QN => n4696);
   registers_reg_10_20_inst : DFF_X1 port map( D => n7875, CK => clk, Q => 
                           n10267, QN => n4697);
   registers_reg_10_19_inst : DFF_X1 port map( D => n7874, CK => clk, Q => 
                           n10335, QN => n4698);
   registers_reg_10_18_inst : DFF_X1 port map( D => n7873, CK => clk, Q => 
                           n10402, QN => n4699);
   registers_reg_10_17_inst : DFF_X1 port map( D => n7872, CK => clk, Q => 
                           n10469, QN => n4700);
   registers_reg_10_16_inst : DFF_X1 port map( D => n7871, CK => clk, Q => 
                           n10537, QN => n4701);
   registers_reg_10_15_inst : DFF_X1 port map( D => n7870, CK => clk, Q => 
                           n10604, QN => n4702);
   registers_reg_10_14_inst : DFF_X1 port map( D => n7869, CK => clk, Q => 
                           n10671, QN => n4703);
   registers_reg_10_13_inst : DFF_X1 port map( D => n7868, CK => clk, Q => 
                           n10738, QN => n4704);
   registers_reg_10_12_inst : DFF_X1 port map( D => n7867, CK => clk, Q => 
                           n10806, QN => n4705);
   registers_reg_10_11_inst : DFF_X1 port map( D => n7866, CK => clk, Q => 
                           n10873, QN => n4706);
   registers_reg_10_10_inst : DFF_X1 port map( D => n7865, CK => clk, Q => 
                           n10940, QN => n4707);
   registers_reg_10_9_inst : DFF_X1 port map( D => n7864, CK => clk, Q => 
                           n11007, QN => n4708);
   registers_reg_10_8_inst : DFF_X1 port map( D => n7863, CK => clk, Q => 
                           n11075, QN => n4709);
   registers_reg_10_7_inst : DFF_X1 port map( D => n7862, CK => clk, Q => 
                           n11142, QN => n4710);
   registers_reg_10_6_inst : DFF_X1 port map( D => n7861, CK => clk, Q => 
                           n11209, QN => n4711);
   registers_reg_10_5_inst : DFF_X1 port map( D => n7860, CK => clk, Q => 
                           n11276, QN => n4712);
   registers_reg_10_4_inst : DFF_X1 port map( D => n7859, CK => clk, Q => 
                           n11344, QN => n4713);
   registers_reg_9_63_inst : DFF_X1 port map( D => n7854, CK => clk, Q => n3020
                           , QN => n4720);
   registers_reg_9_62_inst : DFF_X1 port map( D => n7853, CK => clk, Q => n3260
                           , QN => n4721);
   registers_reg_9_61_inst : DFF_X1 port map( D => n7852, CK => clk, Q => n4176
                           , QN => n4722);
   registers_reg_9_60_inst : DFF_X1 port map( D => n7851, CK => clk, Q => n5301
                           , QN => n4723);
   registers_reg_9_59_inst : DFF_X1 port map( D => n7850, CK => clk, Q => n5371
                           , QN => n4724);
   registers_reg_9_58_inst : DFF_X1 port map( D => n7849, CK => clk, Q => n5439
                           , QN => n4725);
   registers_reg_9_57_inst : DFF_X1 port map( D => n7848, CK => clk, Q => n5508
                           , QN => n4726);
   registers_reg_9_56_inst : DFF_X1 port map( D => n7847, CK => clk, Q => n5577
                           , QN => n4727);
   registers_reg_9_55_inst : DFF_X1 port map( D => n7846, CK => clk, Q => n5645
                           , QN => n4728);
   registers_reg_9_54_inst : DFF_X1 port map( D => n7845, CK => clk, Q => n5715
                           , QN => n4729);
   registers_reg_9_53_inst : DFF_X1 port map( D => n7844, CK => clk, Q => n5787
                           , QN => n4730);
   registers_reg_9_52_inst : DFF_X1 port map( D => n7843, CK => clk, Q => n5854
                           , QN => n4731);
   registers_reg_9_51_inst : DFF_X1 port map( D => n7842, CK => clk, Q => n5921
                           , QN => n4732);
   registers_reg_9_50_inst : DFF_X1 port map( D => n7841, CK => clk, Q => n5989
                           , QN => n4733);
   registers_reg_9_49_inst : DFF_X1 port map( D => n7840, CK => clk, Q => n6057
                           , QN => n4734);
   registers_reg_9_48_inst : DFF_X1 port map( D => n7839, CK => clk, Q => n6123
                           , QN => n4735);
   registers_reg_9_47_inst : DFF_X1 port map( D => n7838, CK => clk, Q => n6189
                           , QN => n4736);
   registers_reg_9_46_inst : DFF_X1 port map( D => n7837, CK => clk, Q => n6255
                           , QN => n4737);
   registers_reg_9_45_inst : DFF_X1 port map( D => n7836, CK => clk, Q => n6321
                           , QN => n4738);
   registers_reg_9_44_inst : DFF_X1 port map( D => n7835, CK => clk, Q => n6387
                           , QN => n4739);
   registers_reg_9_43_inst : DFF_X1 port map( D => n7834, CK => clk, Q => n6453
                           , QN => n4740);
   registers_reg_9_42_inst : DFF_X1 port map( D => n7833, CK => clk, Q => n6519
                           , QN => n4741);
   registers_reg_9_41_inst : DFF_X1 port map( D => n7832, CK => clk, Q => n6585
                           , QN => n4742);
   registers_reg_9_40_inst : DFF_X1 port map( D => n7831, CK => clk, Q => n6652
                           , QN => n4743);
   registers_reg_9_39_inst : DFF_X1 port map( D => n7830, CK => clk, Q => n6719
                           , QN => n4744);
   registers_reg_9_38_inst : DFF_X1 port map( D => n7829, CK => clk, Q => n6786
                           , QN => n4745);
   registers_reg_9_37_inst : DFF_X1 port map( D => n7828, CK => clk, Q => n6853
                           , QN => n4746);
   registers_reg_9_36_inst : DFF_X1 port map( D => n7827, CK => clk, Q => n6920
                           , QN => n4747);
   registers_reg_9_35_inst : DFF_X1 port map( D => n7826, CK => clk, Q => n6987
                           , QN => n4748);
   registers_reg_9_34_inst : DFF_X1 port map( D => n7825, CK => clk, Q => n9294
                           , QN => n4749);
   registers_reg_9_33_inst : DFF_X1 port map( D => n7824, CK => clk, Q => n9361
                           , QN => n4750);
   registers_reg_9_32_inst : DFF_X1 port map( D => n7823, CK => clk, Q => n9429
                           , QN => n4751);
   registers_reg_9_31_inst : DFF_X1 port map( D => n7822, CK => clk, Q => n9496
                           , QN => n4752);
   registers_reg_9_30_inst : DFF_X1 port map( D => n7821, CK => clk, Q => n9563
                           , QN => n4753);
   registers_reg_9_29_inst : DFF_X1 port map( D => n7820, CK => clk, Q => n9630
                           , QN => n4754);
   registers_reg_9_28_inst : DFF_X1 port map( D => n7819, CK => clk, Q => n9698
                           , QN => n4755);
   registers_reg_9_27_inst : DFF_X1 port map( D => n7818, CK => clk, Q => n9765
                           , QN => n4756);
   registers_reg_9_26_inst : DFF_X1 port map( D => n7817, CK => clk, Q => n9832
                           , QN => n4757);
   registers_reg_9_25_inst : DFF_X1 port map( D => n7816, CK => clk, Q => n9899
                           , QN => n4758);
   registers_reg_9_24_inst : DFF_X1 port map( D => n7815, CK => clk, Q => n9967
                           , QN => n4759);
   registers_reg_9_23_inst : DFF_X1 port map( D => n7814, CK => clk, Q => 
                           n10034, QN => n4760);
   registers_reg_9_22_inst : DFF_X1 port map( D => n7813, CK => clk, Q => 
                           n10101, QN => n4761);
   registers_reg_9_21_inst : DFF_X1 port map( D => n7812, CK => clk, Q => 
                           n10169, QN => n4762);
   registers_reg_9_20_inst : DFF_X1 port map( D => n7811, CK => clk, Q => 
                           n10236, QN => n4763);
   registers_reg_9_19_inst : DFF_X1 port map( D => n7810, CK => clk, Q => 
                           n10303, QN => n4764);
   registers_reg_9_18_inst : DFF_X1 port map( D => n7809, CK => clk, Q => 
                           n10370, QN => n4765);
   registers_reg_9_17_inst : DFF_X1 port map( D => n7808, CK => clk, Q => 
                           n10438, QN => n4766);
   registers_reg_9_16_inst : DFF_X1 port map( D => n7807, CK => clk, Q => 
                           n10505, QN => n4767);
   registers_reg_9_15_inst : DFF_X1 port map( D => n7806, CK => clk, Q => 
                           n10572, QN => n4768);
   registers_reg_9_14_inst : DFF_X1 port map( D => n7805, CK => clk, Q => 
                           n10639, QN => n4769);
   registers_reg_9_13_inst : DFF_X1 port map( D => n7804, CK => clk, Q => 
                           n10707, QN => n4770);
   registers_reg_9_12_inst : DFF_X1 port map( D => n7803, CK => clk, Q => 
                           n10774, QN => n4771);
   registers_reg_9_11_inst : DFF_X1 port map( D => n7802, CK => clk, Q => 
                           n10841, QN => n4772);
   registers_reg_9_10_inst : DFF_X1 port map( D => n7801, CK => clk, Q => 
                           n10909, QN => n4773);
   registers_reg_9_9_inst : DFF_X1 port map( D => n7800, CK => clk, Q => n10976
                           , QN => n4774);
   registers_reg_9_8_inst : DFF_X1 port map( D => n7799, CK => clk, Q => n11043
                           , QN => n4775);
   registers_reg_9_7_inst : DFF_X1 port map( D => n7798, CK => clk, Q => n11110
                           , QN => n4776);
   registers_reg_9_6_inst : DFF_X1 port map( D => n7797, CK => clk, Q => n11178
                           , QN => n4777);
   registers_reg_9_5_inst : DFF_X1 port map( D => n7796, CK => clk, Q => n11245
                           , QN => n4778);
   registers_reg_9_4_inst : DFF_X1 port map( D => n7795, CK => clk, Q => n11312
                           , QN => n4779);
   registers_reg_8_63_inst : DFF_X1 port map( D => n7790, CK => clk, Q => n3192
                           , QN => n4787);
   registers_reg_8_62_inst : DFF_X1 port map( D => n7789, CK => clk, Q => n3571
                           , QN => n4788);
   registers_reg_8_61_inst : DFF_X1 port map( D => n7788, CK => clk, Q => n4853
                           , QN => n4789);
   registers_reg_8_60_inst : DFF_X1 port map( D => n7787, CK => clk, Q => n5338
                           , QN => n4790);
   registers_reg_8_59_inst : DFF_X1 port map( D => n7786, CK => clk, Q => n5408
                           , QN => n4791);
   registers_reg_8_58_inst : DFF_X1 port map( D => n7785, CK => clk, Q => n5476
                           , QN => n4792);
   registers_reg_8_57_inst : DFF_X1 port map( D => n7784, CK => clk, Q => n5545
                           , QN => n4793);
   registers_reg_8_56_inst : DFF_X1 port map( D => n7783, CK => clk, Q => n5614
                           , QN => n4794);
   registers_reg_8_55_inst : DFF_X1 port map( D => n7782, CK => clk, Q => n5682
                           , QN => n4795);
   registers_reg_8_54_inst : DFF_X1 port map( D => n7781, CK => clk, Q => n5752
                           , QN => n4796);
   registers_reg_8_53_inst : DFF_X1 port map( D => n7780, CK => clk, Q => n5824
                           , QN => n4797);
   registers_reg_8_52_inst : DFF_X1 port map( D => n7779, CK => clk, Q => n5891
                           , QN => n4798);
   registers_reg_8_51_inst : DFF_X1 port map( D => n7778, CK => clk, Q => n5958
                           , QN => n4799);
   registers_reg_8_50_inst : DFF_X1 port map( D => n7777, CK => clk, Q => n6026
                           , QN => n4800);
   registers_reg_8_49_inst : DFF_X1 port map( D => n7776, CK => clk, Q => n6094
                           , QN => n4801);
   registers_reg_8_48_inst : DFF_X1 port map( D => n7775, CK => clk, Q => n6160
                           , QN => n4802);
   registers_reg_8_47_inst : DFF_X1 port map( D => n7774, CK => clk, Q => n6226
                           , QN => n4803);
   registers_reg_8_46_inst : DFF_X1 port map( D => n7773, CK => clk, Q => n6292
                           , QN => n4804);
   registers_reg_8_45_inst : DFF_X1 port map( D => n7772, CK => clk, Q => n6358
                           , QN => n4805);
   registers_reg_8_44_inst : DFF_X1 port map( D => n7771, CK => clk, Q => n6424
                           , QN => n4806);
   registers_reg_8_43_inst : DFF_X1 port map( D => n7770, CK => clk, Q => n6490
                           , QN => n4807);
   registers_reg_8_42_inst : DFF_X1 port map( D => n7769, CK => clk, Q => n6556
                           , QN => n4808);
   registers_reg_8_41_inst : DFF_X1 port map( D => n7768, CK => clk, Q => n6622
                           , QN => n4809);
   registers_reg_8_40_inst : DFF_X1 port map( D => n7767, CK => clk, Q => n6689
                           , QN => n4810);
   registers_reg_8_39_inst : DFF_X1 port map( D => n7766, CK => clk, Q => n6757
                           , QN => n4811);
   registers_reg_8_38_inst : DFF_X1 port map( D => n7765, CK => clk, Q => n6824
                           , QN => n4812);
   registers_reg_8_37_inst : DFF_X1 port map( D => n7764, CK => clk, Q => n6891
                           , QN => n4813);
   registers_reg_8_36_inst : DFF_X1 port map( D => n7763, CK => clk, Q => n6958
                           , QN => n4814);
   registers_reg_8_35_inst : DFF_X1 port map( D => n7762, CK => clk, Q => n9264
                           , QN => n4815);
   registers_reg_8_34_inst : DFF_X1 port map( D => n7761, CK => clk, Q => n9332
                           , QN => n4816);
   registers_reg_8_33_inst : DFF_X1 port map( D => n7760, CK => clk, Q => n9399
                           , QN => n4817);
   registers_reg_8_32_inst : DFF_X1 port map( D => n7759, CK => clk, Q => n9466
                           , QN => n4818);
   registers_reg_8_31_inst : DFF_X1 port map( D => n7758, CK => clk, Q => n9534
                           , QN => n4819);
   registers_reg_8_30_inst : DFF_X1 port map( D => n7757, CK => clk, Q => n9601
                           , QN => n4820);
   registers_reg_8_29_inst : DFF_X1 port map( D => n7756, CK => clk, Q => n9668
                           , QN => n4821);
   registers_reg_8_28_inst : DFF_X1 port map( D => n7755, CK => clk, Q => n9735
                           , QN => n4822);
   registers_reg_8_27_inst : DFF_X1 port map( D => n7754, CK => clk, Q => n9803
                           , QN => n4823);
   registers_reg_8_26_inst : DFF_X1 port map( D => n7753, CK => clk, Q => n9870
                           , QN => n4824);
   registers_reg_8_25_inst : DFF_X1 port map( D => n7752, CK => clk, Q => n9937
                           , QN => n4825);
   registers_reg_8_24_inst : DFF_X1 port map( D => n7751, CK => clk, Q => 
                           n10004, QN => n4826);
   registers_reg_8_23_inst : DFF_X1 port map( D => n7750, CK => clk, Q => 
                           n10072, QN => n4827);
   registers_reg_8_22_inst : DFF_X1 port map( D => n7749, CK => clk, Q => 
                           n10139, QN => n4828);
   registers_reg_8_21_inst : DFF_X1 port map( D => n7748, CK => clk, Q => 
                           n10206, QN => n4829);
   registers_reg_8_20_inst : DFF_X1 port map( D => n7747, CK => clk, Q => 
                           n10274, QN => n4830);
   registers_reg_8_19_inst : DFF_X1 port map( D => n7746, CK => clk, Q => 
                           n10341, QN => n4831);
   registers_reg_8_18_inst : DFF_X1 port map( D => n7745, CK => clk, Q => 
                           n10408, QN => n4832);
   registers_reg_8_17_inst : DFF_X1 port map( D => n7744, CK => clk, Q => 
                           n10475, QN => n4833);
   registers_reg_8_16_inst : DFF_X1 port map( D => n7743, CK => clk, Q => 
                           n10543, QN => n4834);
   registers_reg_8_15_inst : DFF_X1 port map( D => n7742, CK => clk, Q => 
                           n10610, QN => n4835);
   registers_reg_8_14_inst : DFF_X1 port map( D => n7741, CK => clk, Q => 
                           n10677, QN => n4836);
   registers_reg_8_13_inst : DFF_X1 port map( D => n7740, CK => clk, Q => 
                           n10744, QN => n4837);
   registers_reg_8_12_inst : DFF_X1 port map( D => n7739, CK => clk, Q => 
                           n10812, QN => n4838);
   registers_reg_8_11_inst : DFF_X1 port map( D => n7738, CK => clk, Q => 
                           n10879, QN => n4839);
   registers_reg_8_10_inst : DFF_X1 port map( D => n7737, CK => clk, Q => 
                           n10946, QN => n4840);
   registers_reg_8_9_inst : DFF_X1 port map( D => n7736, CK => clk, Q => n11014
                           , QN => n4841);
   registers_reg_8_8_inst : DFF_X1 port map( D => n7735, CK => clk, Q => n11081
                           , QN => n4842);
   registers_reg_8_7_inst : DFF_X1 port map( D => n7734, CK => clk, Q => n11148
                           , QN => n4843);
   registers_reg_8_6_inst : DFF_X1 port map( D => n7733, CK => clk, Q => n11215
                           , QN => n4844);
   registers_reg_8_5_inst : DFF_X1 port map( D => n7732, CK => clk, Q => n11283
                           , QN => n4845);
   registers_reg_8_4_inst : DFF_X1 port map( D => n7731, CK => clk, Q => n11350
                           , QN => n4846);
   registers_reg_30_63_inst : DFF_X1 port map( D => n9198, CK => clk, Q => 
                           n18689, QN => n3303);
   registers_reg_30_62_inst : DFF_X1 port map( D => n9197, CK => clk, Q => 
                           n18688, QN => n3304);
   registers_reg_30_61_inst : DFF_X1 port map( D => n9196, CK => clk, Q => 
                           n18687, QN => n3305);
   registers_reg_30_60_inst : DFF_X1 port map( D => n9195, CK => clk, Q => 
                           n18686, QN => n3306);
   registers_reg_30_59_inst : DFF_X1 port map( D => n9194, CK => clk, Q => 
                           n18685, QN => n3307);
   registers_reg_30_58_inst : DFF_X1 port map( D => n9193, CK => clk, Q => 
                           n18684, QN => n3308);
   registers_reg_30_57_inst : DFF_X1 port map( D => n9192, CK => clk, Q => 
                           n18683, QN => n3309);
   registers_reg_30_56_inst : DFF_X1 port map( D => n9191, CK => clk, Q => 
                           n18682, QN => n3310);
   registers_reg_30_55_inst : DFF_X1 port map( D => n9190, CK => clk, Q => 
                           n18681, QN => n3311);
   registers_reg_15_3_inst : DFF_X1 port map( D => n8178, CK => clk, Q => 
                           registers_15_3_port, QN => n2010);
   registers_reg_15_2_inst : DFF_X1 port map( D => n8177, CK => clk, Q => 
                           registers_15_2_port, QN => n2011);
   registers_reg_15_1_inst : DFF_X1 port map( D => n8176, CK => clk, Q => 
                           registers_15_1_port, QN => n2012);
   registers_reg_15_0_inst : DFF_X1 port map( D => n8175, CK => clk, Q => 
                           registers_15_0_port, QN => n2013);
   registers_reg_14_3_inst : DFF_X1 port map( D => n8114, CK => clk, Q => 
                           registers_14_3_port, QN => n2078);
   registers_reg_14_2_inst : DFF_X1 port map( D => n8113, CK => clk, Q => 
                           registers_14_2_port, QN => n2079);
   registers_reg_14_1_inst : DFF_X1 port map( D => n8112, CK => clk, Q => 
                           registers_14_1_port, QN => n2080);
   registers_reg_14_0_inst : DFF_X1 port map( D => n8111, CK => clk, Q => 
                           registers_14_0_port, QN => n2081);
   registers_reg_11_3_inst : DFF_X1 port map( D => n7922, CK => clk, Q => 
                           n18680, QN => n2183);
   registers_reg_11_2_inst : DFF_X1 port map( D => n7921, CK => clk, Q => 
                           n18679, QN => n2186);
   registers_reg_11_1_inst : DFF_X1 port map( D => n7920, CK => clk, Q => 
                           n18678, QN => n2189);
   registers_reg_11_0_inst : DFF_X1 port map( D => n7919, CK => clk, Q => 
                           n18677, QN => n2192);
   registers_reg_2_3_inst : DFF_X1 port map( D => n7346, CK => clk, Q => n18676
                           , QN => n2760);
   registers_reg_2_2_inst : DFF_X1 port map( D => n7345, CK => clk, Q => n18675
                           , QN => n2761);
   registers_reg_2_1_inst : DFF_X1 port map( D => n7344, CK => clk, Q => n18674
                           , QN => n2762);
   registers_reg_2_0_inst : DFF_X1 port map( D => n7343, CK => clk, Q => n18673
                           , QN => n2763);
   registers_reg_3_3_inst : DFF_X1 port map( D => n7410, CK => clk, Q => 
                           registers_3_3_port, QN => n2438);
   registers_reg_3_2_inst : DFF_X1 port map( D => n7409, CK => clk, Q => 
                           registers_3_2_port, QN => n2439);
   registers_reg_3_1_inst : DFF_X1 port map( D => n7408, CK => clk, Q => 
                           registers_3_1_port, QN => n2440);
   registers_reg_3_0_inst : DFF_X1 port map( D => n7407, CK => clk, Q => 
                           registers_3_0_port, QN => n2441);
   registers_reg_0_63_inst : DFF_X1 port map( D => n7278, CK => clk, Q => 
                           n18672, QN => n2768);
   registers_reg_0_62_inst : DFF_X1 port map( D => n7274, CK => clk, Q => 
                           n18671, QN => n3208);
   registers_reg_0_61_inst : DFF_X1 port map( D => n7270, CK => clk, Q => 
                           n18670, QN => n3638);
   registers_reg_0_60_inst : DFF_X1 port map( D => n7266, CK => clk, Q => 
                           n18669, QN => n4856);
   registers_reg_18_3_inst : DFF_X1 port map( D => n8370, CK => clk, Q => 
                           n18668, QN => n1934);
   registers_reg_18_2_inst : DFF_X1 port map( D => n8369, CK => clk, Q => 
                           n18667, QN => n1935);
   registers_reg_18_1_inst : DFF_X1 port map( D => n8368, CK => clk, Q => 
                           n18666, QN => n1936);
   registers_reg_18_0_inst : DFF_X1 port map( D => n8367, CK => clk, Q => 
                           n18665, QN => n1937);
   registers_reg_14_63_inst : DFF_X1 port map( D => n8174, CK => clk, Q => 
                           registers_14_63_port, QN => n2018);
   registers_reg_14_62_inst : DFF_X1 port map( D => n8173, CK => clk, Q => 
                           registers_14_62_port, QN => n2019);
   registers_reg_14_61_inst : DFF_X1 port map( D => n8172, CK => clk, Q => 
                           registers_14_61_port, QN => n2020);
   registers_reg_14_60_inst : DFF_X1 port map( D => n8171, CK => clk, Q => 
                           registers_14_60_port, QN => n2021);
   registers_reg_14_59_inst : DFF_X1 port map( D => n8170, CK => clk, Q => 
                           registers_14_59_port, QN => n2022);
   registers_reg_14_58_inst : DFF_X1 port map( D => n8169, CK => clk, Q => 
                           registers_14_58_port, QN => n2023);
   registers_reg_14_57_inst : DFF_X1 port map( D => n8168, CK => clk, Q => 
                           registers_14_57_port, QN => n2024);
   registers_reg_14_56_inst : DFF_X1 port map( D => n8167, CK => clk, Q => 
                           registers_14_56_port, QN => n2025);
   registers_reg_14_55_inst : DFF_X1 port map( D => n8166, CK => clk, Q => 
                           registers_14_55_port, QN => n2026);
   registers_reg_14_54_inst : DFF_X1 port map( D => n8165, CK => clk, Q => 
                           registers_14_54_port, QN => n2027);
   registers_reg_14_53_inst : DFF_X1 port map( D => n8164, CK => clk, Q => 
                           registers_14_53_port, QN => n2028);
   registers_reg_14_52_inst : DFF_X1 port map( D => n8163, CK => clk, Q => 
                           registers_14_52_port, QN => n2029);
   registers_reg_14_51_inst : DFF_X1 port map( D => n8162, CK => clk, Q => 
                           registers_14_51_port, QN => n2030);
   registers_reg_14_50_inst : DFF_X1 port map( D => n8161, CK => clk, Q => 
                           registers_14_50_port, QN => n2031);
   registers_reg_14_49_inst : DFF_X1 port map( D => n8160, CK => clk, Q => 
                           registers_14_49_port, QN => n2032);
   registers_reg_14_48_inst : DFF_X1 port map( D => n8159, CK => clk, Q => 
                           registers_14_48_port, QN => n2033);
   registers_reg_14_47_inst : DFF_X1 port map( D => n8158, CK => clk, Q => 
                           registers_14_47_port, QN => n2034);
   registers_reg_14_46_inst : DFF_X1 port map( D => n8157, CK => clk, Q => 
                           registers_14_46_port, QN => n2035);
   registers_reg_14_45_inst : DFF_X1 port map( D => n8156, CK => clk, Q => 
                           registers_14_45_port, QN => n2036);
   registers_reg_14_44_inst : DFF_X1 port map( D => n8155, CK => clk, Q => 
                           registers_14_44_port, QN => n2037);
   registers_reg_14_43_inst : DFF_X1 port map( D => n8154, CK => clk, Q => 
                           registers_14_43_port, QN => n2038);
   registers_reg_14_42_inst : DFF_X1 port map( D => n8153, CK => clk, Q => 
                           registers_14_42_port, QN => n2039);
   registers_reg_14_41_inst : DFF_X1 port map( D => n8152, CK => clk, Q => 
                           registers_14_41_port, QN => n2040);
   registers_reg_14_40_inst : DFF_X1 port map( D => n8151, CK => clk, Q => 
                           registers_14_40_port, QN => n2041);
   registers_reg_14_39_inst : DFF_X1 port map( D => n8150, CK => clk, Q => 
                           registers_14_39_port, QN => n2042);
   registers_reg_14_38_inst : DFF_X1 port map( D => n8149, CK => clk, Q => 
                           registers_14_38_port, QN => n2043);
   registers_reg_14_37_inst : DFF_X1 port map( D => n8148, CK => clk, Q => 
                           registers_14_37_port, QN => n2044);
   registers_reg_14_36_inst : DFF_X1 port map( D => n8147, CK => clk, Q => 
                           registers_14_36_port, QN => n2045);
   registers_reg_14_35_inst : DFF_X1 port map( D => n8146, CK => clk, Q => 
                           registers_14_35_port, QN => n2046);
   registers_reg_14_34_inst : DFF_X1 port map( D => n8145, CK => clk, Q => 
                           registers_14_34_port, QN => n2047);
   registers_reg_14_33_inst : DFF_X1 port map( D => n8144, CK => clk, Q => 
                           registers_14_33_port, QN => n2048);
   registers_reg_14_32_inst : DFF_X1 port map( D => n8143, CK => clk, Q => 
                           registers_14_32_port, QN => n2049);
   registers_reg_14_31_inst : DFF_X1 port map( D => n8142, CK => clk, Q => 
                           registers_14_31_port, QN => n2050);
   registers_reg_14_30_inst : DFF_X1 port map( D => n8141, CK => clk, Q => 
                           registers_14_30_port, QN => n2051);
   registers_reg_14_29_inst : DFF_X1 port map( D => n8140, CK => clk, Q => 
                           registers_14_29_port, QN => n2052);
   registers_reg_14_28_inst : DFF_X1 port map( D => n8139, CK => clk, Q => 
                           registers_14_28_port, QN => n2053);
   registers_reg_14_27_inst : DFF_X1 port map( D => n8138, CK => clk, Q => 
                           registers_14_27_port, QN => n2054);
   registers_reg_14_26_inst : DFF_X1 port map( D => n8137, CK => clk, Q => 
                           registers_14_26_port, QN => n2055);
   registers_reg_14_25_inst : DFF_X1 port map( D => n8136, CK => clk, Q => 
                           registers_14_25_port, QN => n2056);
   registers_reg_14_24_inst : DFF_X1 port map( D => n8135, CK => clk, Q => 
                           registers_14_24_port, QN => n2057);
   registers_reg_14_23_inst : DFF_X1 port map( D => n8134, CK => clk, Q => 
                           registers_14_23_port, QN => n2058);
   registers_reg_14_22_inst : DFF_X1 port map( D => n8133, CK => clk, Q => 
                           registers_14_22_port, QN => n2059);
   registers_reg_14_21_inst : DFF_X1 port map( D => n8132, CK => clk, Q => 
                           registers_14_21_port, QN => n2060);
   registers_reg_14_20_inst : DFF_X1 port map( D => n8131, CK => clk, Q => 
                           registers_14_20_port, QN => n2061);
   registers_reg_14_19_inst : DFF_X1 port map( D => n8130, CK => clk, Q => 
                           registers_14_19_port, QN => n2062);
   registers_reg_14_18_inst : DFF_X1 port map( D => n8129, CK => clk, Q => 
                           registers_14_18_port, QN => n2063);
   registers_reg_14_17_inst : DFF_X1 port map( D => n8128, CK => clk, Q => 
                           registers_14_17_port, QN => n2064);
   registers_reg_14_16_inst : DFF_X1 port map( D => n8127, CK => clk, Q => 
                           registers_14_16_port, QN => n2065);
   registers_reg_14_15_inst : DFF_X1 port map( D => n8126, CK => clk, Q => 
                           registers_14_15_port, QN => n2066);
   registers_reg_14_14_inst : DFF_X1 port map( D => n8125, CK => clk, Q => 
                           registers_14_14_port, QN => n2067);
   registers_reg_14_13_inst : DFF_X1 port map( D => n8124, CK => clk, Q => 
                           registers_14_13_port, QN => n2068);
   registers_reg_14_12_inst : DFF_X1 port map( D => n8123, CK => clk, Q => 
                           registers_14_12_port, QN => n2069);
   registers_reg_14_11_inst : DFF_X1 port map( D => n8122, CK => clk, Q => 
                           registers_14_11_port, QN => n2070);
   registers_reg_14_10_inst : DFF_X1 port map( D => n8121, CK => clk, Q => 
                           registers_14_10_port, QN => n2071);
   registers_reg_14_9_inst : DFF_X1 port map( D => n8120, CK => clk, Q => 
                           registers_14_9_port, QN => n2072);
   registers_reg_14_8_inst : DFF_X1 port map( D => n8119, CK => clk, Q => 
                           registers_14_8_port, QN => n2073);
   registers_reg_14_7_inst : DFF_X1 port map( D => n8118, CK => clk, Q => 
                           registers_14_7_port, QN => n2074);
   registers_reg_14_6_inst : DFF_X1 port map( D => n8117, CK => clk, Q => 
                           registers_14_6_port, QN => n2075);
   registers_reg_14_5_inst : DFF_X1 port map( D => n8116, CK => clk, Q => 
                           registers_14_5_port, QN => n2076);
   registers_reg_14_4_inst : DFF_X1 port map( D => n8115, CK => clk, Q => 
                           registers_14_4_port, QN => n2077);
   registers_reg_15_63_inst : DFF_X1 port map( D => n8238, CK => clk, Q => 
                           registers_15_63_port, QN => n1950);
   registers_reg_15_62_inst : DFF_X1 port map( D => n8237, CK => clk, Q => 
                           registers_15_62_port, QN => n1951);
   registers_reg_15_61_inst : DFF_X1 port map( D => n8236, CK => clk, Q => 
                           registers_15_61_port, QN => n1952);
   registers_reg_15_60_inst : DFF_X1 port map( D => n8235, CK => clk, Q => 
                           registers_15_60_port, QN => n1953);
   registers_reg_15_59_inst : DFF_X1 port map( D => n8234, CK => clk, Q => 
                           registers_15_59_port, QN => n1954);
   registers_reg_15_58_inst : DFF_X1 port map( D => n8233, CK => clk, Q => 
                           registers_15_58_port, QN => n1955);
   registers_reg_15_57_inst : DFF_X1 port map( D => n8232, CK => clk, Q => 
                           registers_15_57_port, QN => n1956);
   registers_reg_15_56_inst : DFF_X1 port map( D => n8231, CK => clk, Q => 
                           registers_15_56_port, QN => n1957);
   registers_reg_15_55_inst : DFF_X1 port map( D => n8230, CK => clk, Q => 
                           registers_15_55_port, QN => n1958);
   registers_reg_15_54_inst : DFF_X1 port map( D => n8229, CK => clk, Q => 
                           registers_15_54_port, QN => n1959);
   registers_reg_15_53_inst : DFF_X1 port map( D => n8228, CK => clk, Q => 
                           registers_15_53_port, QN => n1960);
   registers_reg_15_52_inst : DFF_X1 port map( D => n8227, CK => clk, Q => 
                           registers_15_52_port, QN => n1961);
   registers_reg_15_51_inst : DFF_X1 port map( D => n8226, CK => clk, Q => 
                           registers_15_51_port, QN => n1962);
   registers_reg_15_50_inst : DFF_X1 port map( D => n8225, CK => clk, Q => 
                           registers_15_50_port, QN => n1963);
   registers_reg_15_49_inst : DFF_X1 port map( D => n8224, CK => clk, Q => 
                           registers_15_49_port, QN => n1964);
   registers_reg_15_48_inst : DFF_X1 port map( D => n8223, CK => clk, Q => 
                           registers_15_48_port, QN => n1965);
   registers_reg_15_47_inst : DFF_X1 port map( D => n8222, CK => clk, Q => 
                           registers_15_47_port, QN => n1966);
   registers_reg_15_46_inst : DFF_X1 port map( D => n8221, CK => clk, Q => 
                           registers_15_46_port, QN => n1967);
   registers_reg_15_45_inst : DFF_X1 port map( D => n8220, CK => clk, Q => 
                           registers_15_45_port, QN => n1968);
   registers_reg_15_44_inst : DFF_X1 port map( D => n8219, CK => clk, Q => 
                           registers_15_44_port, QN => n1969);
   registers_reg_15_43_inst : DFF_X1 port map( D => n8218, CK => clk, Q => 
                           registers_15_43_port, QN => n1970);
   registers_reg_15_42_inst : DFF_X1 port map( D => n8217, CK => clk, Q => 
                           registers_15_42_port, QN => n1971);
   registers_reg_15_41_inst : DFF_X1 port map( D => n8216, CK => clk, Q => 
                           registers_15_41_port, QN => n1972);
   registers_reg_15_40_inst : DFF_X1 port map( D => n8215, CK => clk, Q => 
                           registers_15_40_port, QN => n1973);
   registers_reg_15_39_inst : DFF_X1 port map( D => n8214, CK => clk, Q => 
                           registers_15_39_port, QN => n1974);
   registers_reg_15_38_inst : DFF_X1 port map( D => n8213, CK => clk, Q => 
                           registers_15_38_port, QN => n1975);
   registers_reg_15_37_inst : DFF_X1 port map( D => n8212, CK => clk, Q => 
                           registers_15_37_port, QN => n1976);
   registers_reg_15_36_inst : DFF_X1 port map( D => n8211, CK => clk, Q => 
                           registers_15_36_port, QN => n1977);
   registers_reg_15_35_inst : DFF_X1 port map( D => n8210, CK => clk, Q => 
                           registers_15_35_port, QN => n1978);
   registers_reg_15_34_inst : DFF_X1 port map( D => n8209, CK => clk, Q => 
                           registers_15_34_port, QN => n1979);
   registers_reg_15_33_inst : DFF_X1 port map( D => n8208, CK => clk, Q => 
                           registers_15_33_port, QN => n1980);
   registers_reg_15_32_inst : DFF_X1 port map( D => n8207, CK => clk, Q => 
                           registers_15_32_port, QN => n1981);
   registers_reg_15_31_inst : DFF_X1 port map( D => n8206, CK => clk, Q => 
                           registers_15_31_port, QN => n1982);
   registers_reg_15_30_inst : DFF_X1 port map( D => n8205, CK => clk, Q => 
                           registers_15_30_port, QN => n1983);
   registers_reg_15_29_inst : DFF_X1 port map( D => n8204, CK => clk, Q => 
                           registers_15_29_port, QN => n1984);
   registers_reg_15_28_inst : DFF_X1 port map( D => n8203, CK => clk, Q => 
                           registers_15_28_port, QN => n1985);
   registers_reg_15_27_inst : DFF_X1 port map( D => n8202, CK => clk, Q => 
                           registers_15_27_port, QN => n1986);
   registers_reg_15_26_inst : DFF_X1 port map( D => n8201, CK => clk, Q => 
                           registers_15_26_port, QN => n1987);
   registers_reg_15_25_inst : DFF_X1 port map( D => n8200, CK => clk, Q => 
                           registers_15_25_port, QN => n1988);
   registers_reg_15_24_inst : DFF_X1 port map( D => n8199, CK => clk, Q => 
                           registers_15_24_port, QN => n1989);
   registers_reg_15_23_inst : DFF_X1 port map( D => n8198, CK => clk, Q => 
                           registers_15_23_port, QN => n1990);
   registers_reg_15_22_inst : DFF_X1 port map( D => n8197, CK => clk, Q => 
                           registers_15_22_port, QN => n1991);
   registers_reg_15_21_inst : DFF_X1 port map( D => n8196, CK => clk, Q => 
                           registers_15_21_port, QN => n1992);
   registers_reg_15_20_inst : DFF_X1 port map( D => n8195, CK => clk, Q => 
                           registers_15_20_port, QN => n1993);
   registers_reg_15_19_inst : DFF_X1 port map( D => n8194, CK => clk, Q => 
                           registers_15_19_port, QN => n1994);
   registers_reg_15_18_inst : DFF_X1 port map( D => n8193, CK => clk, Q => 
                           registers_15_18_port, QN => n1995);
   registers_reg_15_17_inst : DFF_X1 port map( D => n8192, CK => clk, Q => 
                           registers_15_17_port, QN => n1996);
   registers_reg_15_16_inst : DFF_X1 port map( D => n8191, CK => clk, Q => 
                           registers_15_16_port, QN => n1997);
   registers_reg_15_15_inst : DFF_X1 port map( D => n8190, CK => clk, Q => 
                           registers_15_15_port, QN => n1998);
   registers_reg_15_14_inst : DFF_X1 port map( D => n8189, CK => clk, Q => 
                           registers_15_14_port, QN => n1999);
   registers_reg_15_13_inst : DFF_X1 port map( D => n8188, CK => clk, Q => 
                           registers_15_13_port, QN => n2000);
   registers_reg_15_12_inst : DFF_X1 port map( D => n8187, CK => clk, Q => 
                           registers_15_12_port, QN => n2001);
   registers_reg_15_11_inst : DFF_X1 port map( D => n8186, CK => clk, Q => 
                           registers_15_11_port, QN => n2002);
   registers_reg_15_10_inst : DFF_X1 port map( D => n8185, CK => clk, Q => 
                           registers_15_10_port, QN => n2003);
   registers_reg_15_9_inst : DFF_X1 port map( D => n8184, CK => clk, Q => 
                           registers_15_9_port, QN => n2004);
   registers_reg_15_8_inst : DFF_X1 port map( D => n8183, CK => clk, Q => 
                           registers_15_8_port, QN => n2005);
   registers_reg_15_7_inst : DFF_X1 port map( D => n8182, CK => clk, Q => 
                           registers_15_7_port, QN => n2006);
   registers_reg_15_6_inst : DFF_X1 port map( D => n8181, CK => clk, Q => 
                           registers_15_6_port, QN => n2007);
   registers_reg_15_5_inst : DFF_X1 port map( D => n8180, CK => clk, Q => 
                           registers_15_5_port, QN => n2008);
   registers_reg_15_4_inst : DFF_X1 port map( D => n8179, CK => clk, Q => 
                           registers_15_4_port, QN => n2009);
   registers_reg_4_3_inst : DFF_X1 port map( D => n7474, CK => clk, Q => 
                           registers_4_3_port, QN => n2371);
   registers_reg_4_2_inst : DFF_X1 port map( D => n7473, CK => clk, Q => 
                           registers_4_2_port, QN => n2372);
   registers_reg_4_1_inst : DFF_X1 port map( D => n7472, CK => clk, Q => 
                           registers_4_1_port, QN => n2373);
   registers_reg_4_0_inst : DFF_X1 port map( D => n7471, CK => clk, Q => 
                           registers_4_0_port, QN => n2374);
   registers_reg_22_3_inst : DFF_X1 port map( D => n8626, CK => clk, Q => 
                           n18664, QN => n1793);
   registers_reg_22_2_inst : DFF_X1 port map( D => n8625, CK => clk, Q => 
                           n18663, QN => n1794);
   registers_reg_22_1_inst : DFF_X1 port map( D => n8624, CK => clk, Q => 
                           n18662, QN => n1795);
   registers_reg_22_0_inst : DFF_X1 port map( D => n8623, CK => clk, Q => 
                           n18661, QN => n1796);
   registers_reg_2_63_inst : DFF_X1 port map( D => n7406, CK => clk, Q => 
                           n18660, QN => n2444);
   registers_reg_2_62_inst : DFF_X1 port map( D => n7405, CK => clk, Q => 
                           n18659, QN => n2445);
   registers_reg_2_61_inst : DFF_X1 port map( D => n7404, CK => clk, Q => 
                           n18658, QN => n2446);
   registers_reg_2_60_inst : DFF_X1 port map( D => n7403, CK => clk, Q => 
                           n18657, QN => n2447);
   registers_reg_2_59_inst : DFF_X1 port map( D => n7402, CK => clk, Q => 
                           n18656, QN => n2448);
   registers_reg_2_58_inst : DFF_X1 port map( D => n7401, CK => clk, Q => 
                           n18655, QN => n2449);
   registers_reg_2_57_inst : DFF_X1 port map( D => n7400, CK => clk, Q => 
                           n18654, QN => n2450);
   registers_reg_2_56_inst : DFF_X1 port map( D => n7399, CK => clk, Q => 
                           n18653, QN => n2451);
   registers_reg_2_55_inst : DFF_X1 port map( D => n7398, CK => clk, Q => 
                           n18652, QN => n2452);
   registers_reg_2_54_inst : DFF_X1 port map( D => n7397, CK => clk, Q => 
                           n18651, QN => n2453);
   registers_reg_2_53_inst : DFF_X1 port map( D => n7396, CK => clk, Q => 
                           n18650, QN => n2454);
   registers_reg_2_52_inst : DFF_X1 port map( D => n7395, CK => clk, Q => 
                           n18649, QN => n2455);
   registers_reg_2_51_inst : DFF_X1 port map( D => n7394, CK => clk, Q => 
                           n18648, QN => n2456);
   registers_reg_2_50_inst : DFF_X1 port map( D => n7393, CK => clk, Q => 
                           n18647, QN => n2457);
   registers_reg_2_49_inst : DFF_X1 port map( D => n7392, CK => clk, Q => 
                           n18646, QN => n2458);
   registers_reg_2_48_inst : DFF_X1 port map( D => n7391, CK => clk, Q => 
                           n18645, QN => n2459);
   registers_reg_2_47_inst : DFF_X1 port map( D => n7390, CK => clk, Q => 
                           n18644, QN => n2460);
   registers_reg_2_46_inst : DFF_X1 port map( D => n7389, CK => clk, Q => 
                           n18643, QN => n2461);
   registers_reg_2_45_inst : DFF_X1 port map( D => n7388, CK => clk, Q => 
                           n18642, QN => n2462);
   registers_reg_2_44_inst : DFF_X1 port map( D => n7387, CK => clk, Q => 
                           n18641, QN => n2463);
   registers_reg_2_43_inst : DFF_X1 port map( D => n7386, CK => clk, Q => 
                           n18640, QN => n2720);
   registers_reg_2_42_inst : DFF_X1 port map( D => n7385, CK => clk, Q => 
                           n18639, QN => n2721);
   registers_reg_2_41_inst : DFF_X1 port map( D => n7384, CK => clk, Q => 
                           n18638, QN => n2722);
   registers_reg_2_40_inst : DFF_X1 port map( D => n7383, CK => clk, Q => 
                           n18637, QN => n2723);
   registers_reg_2_39_inst : DFF_X1 port map( D => n7382, CK => clk, Q => 
                           n18636, QN => n2724);
   registers_reg_2_38_inst : DFF_X1 port map( D => n7381, CK => clk, Q => 
                           n18635, QN => n2725);
   registers_reg_2_37_inst : DFF_X1 port map( D => n7380, CK => clk, Q => 
                           n18634, QN => n2726);
   registers_reg_2_36_inst : DFF_X1 port map( D => n7379, CK => clk, Q => 
                           n18633, QN => n2727);
   registers_reg_2_35_inst : DFF_X1 port map( D => n7378, CK => clk, Q => 
                           n18632, QN => n2728);
   registers_reg_2_34_inst : DFF_X1 port map( D => n7377, CK => clk, Q => 
                           n18631, QN => n2729);
   registers_reg_2_33_inst : DFF_X1 port map( D => n7376, CK => clk, Q => 
                           n18630, QN => n2730);
   registers_reg_2_32_inst : DFF_X1 port map( D => n7375, CK => clk, Q => 
                           n18629, QN => n2731);
   registers_reg_2_31_inst : DFF_X1 port map( D => n7374, CK => clk, Q => 
                           n18628, QN => n2732);
   registers_reg_2_30_inst : DFF_X1 port map( D => n7373, CK => clk, Q => 
                           n18627, QN => n2733);
   registers_reg_2_29_inst : DFF_X1 port map( D => n7372, CK => clk, Q => 
                           n18626, QN => n2734);
   registers_reg_2_28_inst : DFF_X1 port map( D => n7371, CK => clk, Q => 
                           n18625, QN => n2735);
   registers_reg_2_27_inst : DFF_X1 port map( D => n7370, CK => clk, Q => 
                           n18624, QN => n2736);
   registers_reg_2_26_inst : DFF_X1 port map( D => n7369, CK => clk, Q => 
                           n18623, QN => n2737);
   registers_reg_2_25_inst : DFF_X1 port map( D => n7368, CK => clk, Q => 
                           n18622, QN => n2738);
   registers_reg_2_24_inst : DFF_X1 port map( D => n7367, CK => clk, Q => 
                           n18621, QN => n2739);
   registers_reg_2_23_inst : DFF_X1 port map( D => n7366, CK => clk, Q => 
                           n18620, QN => n2740);
   registers_reg_2_22_inst : DFF_X1 port map( D => n7365, CK => clk, Q => 
                           n18619, QN => n2741);
   registers_reg_2_21_inst : DFF_X1 port map( D => n7364, CK => clk, Q => 
                           n18618, QN => n2742);
   registers_reg_2_20_inst : DFF_X1 port map( D => n7363, CK => clk, Q => 
                           n18617, QN => n2743);
   registers_reg_2_19_inst : DFF_X1 port map( D => n7362, CK => clk, Q => 
                           n18616, QN => n2744);
   registers_reg_2_18_inst : DFF_X1 port map( D => n7361, CK => clk, Q => 
                           n18615, QN => n2745);
   registers_reg_2_17_inst : DFF_X1 port map( D => n7360, CK => clk, Q => 
                           n18614, QN => n2746);
   registers_reg_2_16_inst : DFF_X1 port map( D => n7359, CK => clk, Q => 
                           n18613, QN => n2747);
   registers_reg_2_15_inst : DFF_X1 port map( D => n7358, CK => clk, Q => 
                           n18612, QN => n2748);
   registers_reg_2_14_inst : DFF_X1 port map( D => n7357, CK => clk, Q => 
                           n18611, QN => n2749);
   registers_reg_2_13_inst : DFF_X1 port map( D => n7356, CK => clk, Q => 
                           n18610, QN => n2750);
   registers_reg_2_12_inst : DFF_X1 port map( D => n7355, CK => clk, Q => 
                           n18609, QN => n2751);
   registers_reg_2_11_inst : DFF_X1 port map( D => n7354, CK => clk, Q => 
                           n18608, QN => n2752);
   registers_reg_2_10_inst : DFF_X1 port map( D => n7353, CK => clk, Q => 
                           n18607, QN => n2753);
   registers_reg_2_9_inst : DFF_X1 port map( D => n7352, CK => clk, Q => n18606
                           , QN => n2754);
   registers_reg_2_8_inst : DFF_X1 port map( D => n7351, CK => clk, Q => n18605
                           , QN => n2755);
   registers_reg_2_7_inst : DFF_X1 port map( D => n7350, CK => clk, Q => n18604
                           , QN => n2756);
   registers_reg_2_6_inst : DFF_X1 port map( D => n7349, CK => clk, Q => n18603
                           , QN => n2757);
   registers_reg_2_5_inst : DFF_X1 port map( D => n7348, CK => clk, Q => n18602
                           , QN => n2758);
   registers_reg_2_4_inst : DFF_X1 port map( D => n7347, CK => clk, Q => n18601
                           , QN => n2759);
   registers_reg_3_63_inst : DFF_X1 port map( D => n7470, CK => clk, Q => 
                           registers_3_63_port, QN => n2378);
   registers_reg_3_62_inst : DFF_X1 port map( D => n7469, CK => clk, Q => 
                           registers_3_62_port, QN => n2379);
   registers_reg_3_61_inst : DFF_X1 port map( D => n7468, CK => clk, Q => 
                           registers_3_61_port, QN => n2380);
   registers_reg_3_60_inst : DFF_X1 port map( D => n7467, CK => clk, Q => 
                           registers_3_60_port, QN => n2381);
   registers_reg_3_59_inst : DFF_X1 port map( D => n7466, CK => clk, Q => 
                           registers_3_59_port, QN => n2382);
   registers_reg_3_58_inst : DFF_X1 port map( D => n7465, CK => clk, Q => 
                           registers_3_58_port, QN => n2383);
   registers_reg_3_57_inst : DFF_X1 port map( D => n7464, CK => clk, Q => 
                           registers_3_57_port, QN => n2384);
   registers_reg_3_56_inst : DFF_X1 port map( D => n7463, CK => clk, Q => 
                           registers_3_56_port, QN => n2385);
   registers_reg_3_55_inst : DFF_X1 port map( D => n7462, CK => clk, Q => 
                           registers_3_55_port, QN => n2386);
   registers_reg_3_54_inst : DFF_X1 port map( D => n7461, CK => clk, Q => 
                           registers_3_54_port, QN => n2387);
   registers_reg_3_53_inst : DFF_X1 port map( D => n7460, CK => clk, Q => 
                           registers_3_53_port, QN => n2388);
   registers_reg_3_52_inst : DFF_X1 port map( D => n7459, CK => clk, Q => 
                           registers_3_52_port, QN => n2389);
   registers_reg_3_51_inst : DFF_X1 port map( D => n7458, CK => clk, Q => 
                           registers_3_51_port, QN => n2390);
   registers_reg_3_50_inst : DFF_X1 port map( D => n7457, CK => clk, Q => 
                           registers_3_50_port, QN => n2391);
   registers_reg_3_49_inst : DFF_X1 port map( D => n7456, CK => clk, Q => 
                           registers_3_49_port, QN => n2392);
   registers_reg_3_48_inst : DFF_X1 port map( D => n7455, CK => clk, Q => 
                           registers_3_48_port, QN => n2393);
   registers_reg_3_47_inst : DFF_X1 port map( D => n7454, CK => clk, Q => 
                           registers_3_47_port, QN => n2394);
   registers_reg_3_46_inst : DFF_X1 port map( D => n7453, CK => clk, Q => 
                           registers_3_46_port, QN => n2395);
   registers_reg_3_45_inst : DFF_X1 port map( D => n7452, CK => clk, Q => 
                           registers_3_45_port, QN => n2396);
   registers_reg_3_44_inst : DFF_X1 port map( D => n7451, CK => clk, Q => 
                           registers_3_44_port, QN => n2397);
   registers_reg_3_43_inst : DFF_X1 port map( D => n7450, CK => clk, Q => 
                           registers_3_43_port, QN => n2398);
   registers_reg_3_42_inst : DFF_X1 port map( D => n7449, CK => clk, Q => 
                           registers_3_42_port, QN => n2399);
   registers_reg_3_41_inst : DFF_X1 port map( D => n7448, CK => clk, Q => 
                           registers_3_41_port, QN => n2400);
   registers_reg_3_40_inst : DFF_X1 port map( D => n7447, CK => clk, Q => 
                           registers_3_40_port, QN => n2401);
   registers_reg_3_39_inst : DFF_X1 port map( D => n7446, CK => clk, Q => 
                           registers_3_39_port, QN => n2402);
   registers_reg_3_38_inst : DFF_X1 port map( D => n7445, CK => clk, Q => 
                           registers_3_38_port, QN => n2403);
   registers_reg_3_37_inst : DFF_X1 port map( D => n7444, CK => clk, Q => 
                           registers_3_37_port, QN => n2404);
   registers_reg_3_36_inst : DFF_X1 port map( D => n7443, CK => clk, Q => 
                           registers_3_36_port, QN => n2405);
   registers_reg_3_35_inst : DFF_X1 port map( D => n7442, CK => clk, Q => 
                           registers_3_35_port, QN => n2406);
   registers_reg_3_34_inst : DFF_X1 port map( D => n7441, CK => clk, Q => 
                           registers_3_34_port, QN => n2407);
   registers_reg_3_33_inst : DFF_X1 port map( D => n7440, CK => clk, Q => 
                           registers_3_33_port, QN => n2408);
   registers_reg_3_32_inst : DFF_X1 port map( D => n7439, CK => clk, Q => 
                           registers_3_32_port, QN => n2409);
   registers_reg_3_31_inst : DFF_X1 port map( D => n7438, CK => clk, Q => 
                           registers_3_31_port, QN => n2410);
   registers_reg_3_30_inst : DFF_X1 port map( D => n7437, CK => clk, Q => 
                           registers_3_30_port, QN => n2411);
   registers_reg_3_29_inst : DFF_X1 port map( D => n7436, CK => clk, Q => 
                           registers_3_29_port, QN => n2412);
   registers_reg_3_28_inst : DFF_X1 port map( D => n7435, CK => clk, Q => 
                           registers_3_28_port, QN => n2413);
   registers_reg_3_27_inst : DFF_X1 port map( D => n7434, CK => clk, Q => 
                           registers_3_27_port, QN => n2414);
   registers_reg_3_26_inst : DFF_X1 port map( D => n7433, CK => clk, Q => 
                           registers_3_26_port, QN => n2415);
   registers_reg_3_25_inst : DFF_X1 port map( D => n7432, CK => clk, Q => 
                           registers_3_25_port, QN => n2416);
   registers_reg_3_24_inst : DFF_X1 port map( D => n7431, CK => clk, Q => 
                           registers_3_24_port, QN => n2417);
   registers_reg_3_23_inst : DFF_X1 port map( D => n7430, CK => clk, Q => 
                           registers_3_23_port, QN => n2418);
   registers_reg_3_22_inst : DFF_X1 port map( D => n7429, CK => clk, Q => 
                           registers_3_22_port, QN => n2419);
   registers_reg_3_21_inst : DFF_X1 port map( D => n7428, CK => clk, Q => 
                           registers_3_21_port, QN => n2420);
   registers_reg_3_20_inst : DFF_X1 port map( D => n7427, CK => clk, Q => 
                           registers_3_20_port, QN => n2421);
   registers_reg_3_19_inst : DFF_X1 port map( D => n7426, CK => clk, Q => 
                           registers_3_19_port, QN => n2422);
   registers_reg_3_18_inst : DFF_X1 port map( D => n7425, CK => clk, Q => 
                           registers_3_18_port, QN => n2423);
   registers_reg_3_17_inst : DFF_X1 port map( D => n7424, CK => clk, Q => 
                           registers_3_17_port, QN => n2424);
   registers_reg_3_16_inst : DFF_X1 port map( D => n7423, CK => clk, Q => 
                           registers_3_16_port, QN => n2425);
   registers_reg_3_15_inst : DFF_X1 port map( D => n7422, CK => clk, Q => 
                           registers_3_15_port, QN => n2426);
   registers_reg_3_14_inst : DFF_X1 port map( D => n7421, CK => clk, Q => 
                           registers_3_14_port, QN => n2427);
   registers_reg_3_13_inst : DFF_X1 port map( D => n7420, CK => clk, Q => 
                           registers_3_13_port, QN => n2428);
   registers_reg_3_12_inst : DFF_X1 port map( D => n7419, CK => clk, Q => 
                           registers_3_12_port, QN => n2429);
   registers_reg_3_11_inst : DFF_X1 port map( D => n7418, CK => clk, Q => 
                           registers_3_11_port, QN => n2430);
   registers_reg_3_10_inst : DFF_X1 port map( D => n7417, CK => clk, Q => 
                           registers_3_10_port, QN => n2431);
   registers_reg_3_9_inst : DFF_X1 port map( D => n7416, CK => clk, Q => 
                           registers_3_9_port, QN => n2432);
   registers_reg_3_8_inst : DFF_X1 port map( D => n7415, CK => clk, Q => 
                           registers_3_8_port, QN => n2433);
   registers_reg_3_7_inst : DFF_X1 port map( D => n7414, CK => clk, Q => 
                           registers_3_7_port, QN => n2434);
   registers_reg_3_6_inst : DFF_X1 port map( D => n7413, CK => clk, Q => 
                           registers_3_6_port, QN => n2435);
   registers_reg_3_5_inst : DFF_X1 port map( D => n7412, CK => clk, Q => 
                           registers_3_5_port, QN => n2436);
   registers_reg_3_4_inst : DFF_X1 port map( D => n7411, CK => clk, Q => 
                           registers_3_4_port, QN => n2437);
   registers_reg_0_0_inst : DFF_X1 port map( D => n7026, CK => clk, Q => n18600
                           , QN => n11555);
   out_to_mem_reg_63_inst : DFF_X1 port map( D => n7275, CK => clk, Q => 
                           out_to_mem_63_port, QN => n18599);
   out_to_mem_reg_62_inst : DFF_X1 port map( D => n7271, CK => clk, Q => 
                           out_to_mem_62_port, QN => n18598);
   out_to_mem_reg_61_inst : DFF_X1 port map( D => n7267, CK => clk, Q => 
                           out_to_mem_61_port, QN => n18597);
   out_to_mem_reg_60_inst : DFF_X1 port map( D => n7263, CK => clk, Q => 
                           out_to_mem_60_port, QN => n18596);
   registers_reg_21_3_inst : DFF_X1 port map( D => n8562, CK => clk, Q => 
                           n18595, QN => n1860);
   registers_reg_21_2_inst : DFF_X1 port map( D => n8561, CK => clk, Q => 
                           n18594, QN => n1861);
   registers_reg_21_1_inst : DFF_X1 port map( D => n8560, CK => clk, Q => 
                           n18593, QN => n1862);
   registers_reg_21_0_inst : DFF_X1 port map( D => n8559, CK => clk, Q => 
                           n18592, QN => n1863);
   registers_reg_0_11_inst : DFF_X1 port map( D => n7070, CK => clk, Q => 
                           n18591, QN => n10815);
   registers_reg_0_10_inst : DFF_X1 port map( D => n7066, CK => clk, Q => 
                           n18590, QN => n10882);
   registers_reg_0_9_inst : DFF_X1 port map( D => n7062, CK => clk, Q => n18589
                           , QN => n10949);
   registers_reg_0_8_inst : DFF_X1 port map( D => n7058, CK => clk, Q => n18588
                           , QN => n11017);
   registers_reg_0_7_inst : DFF_X1 port map( D => n7054, CK => clk, Q => n18587
                           , QN => n11084);
   registers_reg_0_6_inst : DFF_X1 port map( D => n7050, CK => clk, Q => n18586
                           , QN => n11151);
   registers_reg_0_5_inst : DFF_X1 port map( D => n7046, CK => clk, Q => n18585
                           , QN => n11218);
   registers_reg_0_4_inst : DFF_X1 port map( D => n7042, CK => clk, Q => n18584
                           , QN => n11286);
   registers_reg_0_3_inst : DFF_X1 port map( D => n7038, CK => clk, Q => n18583
                           , QN => n11353);
   registers_reg_0_2_inst : DFF_X1 port map( D => n7034, CK => clk, Q => n18582
                           , QN => n11420);
   registers_reg_0_1_inst : DFF_X1 port map( D => n7030, CK => clk, Q => n18581
                           , QN => n11487);
   registers_reg_0_59_inst : DFF_X1 port map( D => n7262, CK => clk, Q => 
                           n18580, QN => n5341);
   registers_reg_0_58_inst : DFF_X1 port map( D => n7258, CK => clk, Q => 
                           n18579, QN => n5411);
   registers_reg_0_57_inst : DFF_X1 port map( D => n7254, CK => clk, Q => 
                           n18578, QN => n5479);
   registers_reg_0_56_inst : DFF_X1 port map( D => n7250, CK => clk, Q => 
                           n18577, QN => n5548);
   registers_reg_0_55_inst : DFF_X1 port map( D => n7246, CK => clk, Q => 
                           n18576, QN => n5617);
   registers_reg_0_54_inst : DFF_X1 port map( D => n7242, CK => clk, Q => 
                           n18575, QN => n5685);
   registers_reg_0_53_inst : DFF_X1 port map( D => n7238, CK => clk, Q => 
                           n18574, QN => n5755);
   registers_reg_0_52_inst : DFF_X1 port map( D => n7234, CK => clk, Q => 
                           n18573, QN => n5827);
   registers_reg_0_51_inst : DFF_X1 port map( D => n7230, CK => clk, Q => 
                           n18572, QN => n5894);
   registers_reg_0_50_inst : DFF_X1 port map( D => n7226, CK => clk, Q => 
                           n18571, QN => n5961);
   registers_reg_0_49_inst : DFF_X1 port map( D => n7222, CK => clk, Q => 
                           n18570, QN => n6029);
   registers_reg_0_48_inst : DFF_X1 port map( D => n7218, CK => clk, Q => 
                           n18569, QN => n6097);
   registers_reg_0_47_inst : DFF_X1 port map( D => n7214, CK => clk, Q => 
                           n18568, QN => n6163);
   registers_reg_0_46_inst : DFF_X1 port map( D => n7210, CK => clk, Q => 
                           n18567, QN => n6229);
   registers_reg_0_45_inst : DFF_X1 port map( D => n7206, CK => clk, Q => 
                           n18566, QN => n6295);
   registers_reg_0_44_inst : DFF_X1 port map( D => n7202, CK => clk, Q => 
                           n18565, QN => n6361);
   registers_reg_0_43_inst : DFF_X1 port map( D => n7198, CK => clk, Q => 
                           n18564, QN => n6427);
   registers_reg_0_42_inst : DFF_X1 port map( D => n7194, CK => clk, Q => 
                           n18563, QN => n6493);
   registers_reg_0_41_inst : DFF_X1 port map( D => n7190, CK => clk, Q => 
                           n18562, QN => n6559);
   registers_reg_0_40_inst : DFF_X1 port map( D => n7186, CK => clk, Q => 
                           n18561, QN => n6625);
   registers_reg_0_39_inst : DFF_X1 port map( D => n7182, CK => clk, Q => 
                           n18560, QN => n6692);
   registers_reg_0_38_inst : DFF_X1 port map( D => n7178, CK => clk, Q => 
                           n18559, QN => n6760);
   registers_reg_0_37_inst : DFF_X1 port map( D => n7174, CK => clk, Q => 
                           n18558, QN => n6827);
   registers_reg_0_36_inst : DFF_X1 port map( D => n7170, CK => clk, Q => 
                           n18557, QN => n6894);
   registers_reg_0_35_inst : DFF_X1 port map( D => n7166, CK => clk, Q => 
                           n18556, QN => n6961);
   registers_reg_0_34_inst : DFF_X1 port map( D => n7162, CK => clk, Q => 
                           n18555, QN => n9268);
   registers_reg_0_33_inst : DFF_X1 port map( D => n7158, CK => clk, Q => 
                           n18554, QN => n9335);
   registers_reg_0_32_inst : DFF_X1 port map( D => n7154, CK => clk, Q => 
                           n18553, QN => n9402);
   registers_reg_0_31_inst : DFF_X1 port map( D => n7150, CK => clk, Q => 
                           n18552, QN => n9469);
   registers_reg_0_30_inst : DFF_X1 port map( D => n7146, CK => clk, Q => 
                           n18551, QN => n9537);
   registers_reg_0_29_inst : DFF_X1 port map( D => n7142, CK => clk, Q => 
                           n18550, QN => n9604);
   registers_reg_0_28_inst : DFF_X1 port map( D => n7138, CK => clk, Q => 
                           n18549, QN => n9671);
   registers_reg_0_27_inst : DFF_X1 port map( D => n7134, CK => clk, Q => 
                           n18548, QN => n9738);
   registers_reg_0_26_inst : DFF_X1 port map( D => n7130, CK => clk, Q => 
                           n18547, QN => n9806);
   registers_reg_0_25_inst : DFF_X1 port map( D => n7126, CK => clk, Q => 
                           n18546, QN => n9873);
   registers_reg_0_24_inst : DFF_X1 port map( D => n7122, CK => clk, Q => 
                           n18545, QN => n9940);
   registers_reg_0_23_inst : DFF_X1 port map( D => n7118, CK => clk, Q => 
                           n18544, QN => n10008);
   registers_reg_0_22_inst : DFF_X1 port map( D => n7114, CK => clk, Q => 
                           n18543, QN => n10075);
   registers_reg_0_21_inst : DFF_X1 port map( D => n7110, CK => clk, Q => 
                           n18542, QN => n10142);
   registers_reg_0_20_inst : DFF_X1 port map( D => n7106, CK => clk, Q => 
                           n18541, QN => n10209);
   registers_reg_0_19_inst : DFF_X1 port map( D => n7102, CK => clk, Q => 
                           n18540, QN => n10277);
   registers_reg_0_18_inst : DFF_X1 port map( D => n7098, CK => clk, Q => 
                           n18539, QN => n10344);
   registers_reg_0_17_inst : DFF_X1 port map( D => n7094, CK => clk, Q => 
                           n18538, QN => n10411);
   registers_reg_0_16_inst : DFF_X1 port map( D => n7090, CK => clk, Q => 
                           n18537, QN => n10478);
   registers_reg_0_15_inst : DFF_X1 port map( D => n7086, CK => clk, Q => 
                           n18536, QN => n10546);
   registers_reg_0_14_inst : DFF_X1 port map( D => n7082, CK => clk, Q => 
                           n18535, QN => n10613);
   registers_reg_0_13_inst : DFF_X1 port map( D => n7078, CK => clk, Q => 
                           n18534, QN => n10680);
   registers_reg_0_12_inst : DFF_X1 port map( D => n7074, CK => clk, Q => 
                           n18533, QN => n10747);
   registers_reg_18_63_inst : DFF_X1 port map( D => n8430, CK => clk, Q => 
                           n18532, QN => n1874);
   registers_reg_18_62_inst : DFF_X1 port map( D => n8429, CK => clk, Q => 
                           n18531, QN => n1875);
   registers_reg_18_61_inst : DFF_X1 port map( D => n8428, CK => clk, Q => 
                           n18530, QN => n1876);
   registers_reg_18_60_inst : DFF_X1 port map( D => n8427, CK => clk, Q => 
                           n18529, QN => n1877);
   registers_reg_18_59_inst : DFF_X1 port map( D => n8426, CK => clk, Q => 
                           n18528, QN => n1878);
   registers_reg_18_58_inst : DFF_X1 port map( D => n8425, CK => clk, Q => 
                           n18527, QN => n1879);
   registers_reg_18_57_inst : DFF_X1 port map( D => n8424, CK => clk, Q => 
                           n18526, QN => n1880);
   registers_reg_18_56_inst : DFF_X1 port map( D => n8423, CK => clk, Q => 
                           n18525, QN => n1881);
   registers_reg_18_55_inst : DFF_X1 port map( D => n8422, CK => clk, Q => 
                           n18524, QN => n1882);
   registers_reg_18_54_inst : DFF_X1 port map( D => n8421, CK => clk, Q => 
                           n18523, QN => n1883);
   registers_reg_18_53_inst : DFF_X1 port map( D => n8420, CK => clk, Q => 
                           n18522, QN => n1884);
   registers_reg_18_52_inst : DFF_X1 port map( D => n8419, CK => clk, Q => 
                           n18521, QN => n1885);
   registers_reg_18_51_inst : DFF_X1 port map( D => n8418, CK => clk, Q => 
                           n18520, QN => n1886);
   registers_reg_18_50_inst : DFF_X1 port map( D => n8417, CK => clk, Q => 
                           n18519, QN => n1887);
   registers_reg_18_49_inst : DFF_X1 port map( D => n8416, CK => clk, Q => 
                           n18518, QN => n1888);
   registers_reg_18_48_inst : DFF_X1 port map( D => n8415, CK => clk, Q => 
                           n18517, QN => n1889);
   registers_reg_18_47_inst : DFF_X1 port map( D => n8414, CK => clk, Q => 
                           n18516, QN => n1890);
   registers_reg_18_46_inst : DFF_X1 port map( D => n8413, CK => clk, Q => 
                           n18515, QN => n1891);
   registers_reg_18_45_inst : DFF_X1 port map( D => n8412, CK => clk, Q => 
                           n18514, QN => n1892);
   registers_reg_18_44_inst : DFF_X1 port map( D => n8411, CK => clk, Q => 
                           n18513, QN => n1893);
   registers_reg_18_43_inst : DFF_X1 port map( D => n8410, CK => clk, Q => 
                           n18512, QN => n1894);
   registers_reg_18_42_inst : DFF_X1 port map( D => n8409, CK => clk, Q => 
                           n18511, QN => n1895);
   registers_reg_18_41_inst : DFF_X1 port map( D => n8408, CK => clk, Q => 
                           n18510, QN => n1896);
   registers_reg_18_40_inst : DFF_X1 port map( D => n8407, CK => clk, Q => 
                           n18509, QN => n1897);
   registers_reg_18_39_inst : DFF_X1 port map( D => n8406, CK => clk, Q => 
                           n18508, QN => n1898);
   registers_reg_18_38_inst : DFF_X1 port map( D => n8405, CK => clk, Q => 
                           n18507, QN => n1899);
   registers_reg_18_37_inst : DFF_X1 port map( D => n8404, CK => clk, Q => 
                           n18506, QN => n1900);
   registers_reg_18_36_inst : DFF_X1 port map( D => n8403, CK => clk, Q => 
                           n18505, QN => n1901);
   registers_reg_18_35_inst : DFF_X1 port map( D => n8402, CK => clk, Q => 
                           n18504, QN => n1902);
   registers_reg_18_34_inst : DFF_X1 port map( D => n8401, CK => clk, Q => 
                           n18503, QN => n1903);
   registers_reg_18_33_inst : DFF_X1 port map( D => n8400, CK => clk, Q => 
                           n18502, QN => n1904);
   registers_reg_18_32_inst : DFF_X1 port map( D => n8399, CK => clk, Q => 
                           n18501, QN => n1905);
   registers_reg_18_31_inst : DFF_X1 port map( D => n8398, CK => clk, Q => 
                           n18500, QN => n1906);
   registers_reg_18_30_inst : DFF_X1 port map( D => n8397, CK => clk, Q => 
                           n18499, QN => n1907);
   registers_reg_18_29_inst : DFF_X1 port map( D => n8396, CK => clk, Q => 
                           n18498, QN => n1908);
   registers_reg_18_28_inst : DFF_X1 port map( D => n8395, CK => clk, Q => 
                           n18497, QN => n1909);
   registers_reg_18_27_inst : DFF_X1 port map( D => n8394, CK => clk, Q => 
                           n18496, QN => n1910);
   registers_reg_18_26_inst : DFF_X1 port map( D => n8393, CK => clk, Q => 
                           n18495, QN => n1911);
   registers_reg_18_25_inst : DFF_X1 port map( D => n8392, CK => clk, Q => 
                           n18494, QN => n1912);
   registers_reg_18_24_inst : DFF_X1 port map( D => n8391, CK => clk, Q => 
                           n18493, QN => n1913);
   registers_reg_18_23_inst : DFF_X1 port map( D => n8390, CK => clk, Q => 
                           n18492, QN => n1914);
   registers_reg_18_22_inst : DFF_X1 port map( D => n8389, CK => clk, Q => 
                           n18491, QN => n1915);
   registers_reg_18_21_inst : DFF_X1 port map( D => n8388, CK => clk, Q => 
                           n18490, QN => n1916);
   registers_reg_18_20_inst : DFF_X1 port map( D => n8387, CK => clk, Q => 
                           n18489, QN => n1917);
   registers_reg_18_19_inst : DFF_X1 port map( D => n8386, CK => clk, Q => 
                           n18488, QN => n1918);
   registers_reg_18_18_inst : DFF_X1 port map( D => n8385, CK => clk, Q => 
                           n18487, QN => n1919);
   registers_reg_18_17_inst : DFF_X1 port map( D => n8384, CK => clk, Q => 
                           n18486, QN => n1920);
   registers_reg_18_16_inst : DFF_X1 port map( D => n8383, CK => clk, Q => 
                           n18485, QN => n1921);
   registers_reg_18_15_inst : DFF_X1 port map( D => n8382, CK => clk, Q => 
                           n18484, QN => n1922);
   registers_reg_18_14_inst : DFF_X1 port map( D => n8381, CK => clk, Q => 
                           n18483, QN => n1923);
   registers_reg_18_13_inst : DFF_X1 port map( D => n8380, CK => clk, Q => 
                           n18482, QN => n1924);
   registers_reg_18_12_inst : DFF_X1 port map( D => n8379, CK => clk, Q => 
                           n18481, QN => n1925);
   registers_reg_18_11_inst : DFF_X1 port map( D => n8378, CK => clk, Q => 
                           n18480, QN => n1926);
   registers_reg_18_10_inst : DFF_X1 port map( D => n8377, CK => clk, Q => 
                           n18479, QN => n1927);
   registers_reg_18_9_inst : DFF_X1 port map( D => n8376, CK => clk, Q => 
                           n18478, QN => n1928);
   registers_reg_18_8_inst : DFF_X1 port map( D => n8375, CK => clk, Q => 
                           n18477, QN => n1929);
   registers_reg_18_7_inst : DFF_X1 port map( D => n8374, CK => clk, Q => 
                           n18476, QN => n1930);
   registers_reg_18_6_inst : DFF_X1 port map( D => n8373, CK => clk, Q => 
                           n18475, QN => n1931);
   registers_reg_18_5_inst : DFF_X1 port map( D => n8372, CK => clk, Q => 
                           n18474, QN => n1932);
   registers_reg_18_4_inst : DFF_X1 port map( D => n8371, CK => clk, Q => 
                           n18473, QN => n1933);
   registers_reg_11_63_inst : DFF_X1 port map( D => n7982, CK => clk, Q => 
                           n18472, QN => n2097);
   registers_reg_11_62_inst : DFF_X1 port map( D => n7981, CK => clk, Q => 
                           n18471, QN => n2098);
   registers_reg_11_61_inst : DFF_X1 port map( D => n7980, CK => clk, Q => 
                           n18470, QN => n2099);
   registers_reg_11_60_inst : DFF_X1 port map( D => n7979, CK => clk, Q => 
                           n18469, QN => n2100);
   registers_reg_11_59_inst : DFF_X1 port map( D => n7978, CK => clk, Q => 
                           n18468, QN => n2101);
   registers_reg_11_58_inst : DFF_X1 port map( D => n7977, CK => clk, Q => 
                           n18467, QN => n2102);
   registers_reg_11_57_inst : DFF_X1 port map( D => n7976, CK => clk, Q => 
                           n18466, QN => n2103);
   registers_reg_11_56_inst : DFF_X1 port map( D => n7975, CK => clk, Q => 
                           n18465, QN => n2104);
   registers_reg_11_55_inst : DFF_X1 port map( D => n7974, CK => clk, Q => 
                           n18464, QN => n2105);
   registers_reg_11_54_inst : DFF_X1 port map( D => n7973, CK => clk, Q => 
                           n18463, QN => n2106);
   registers_reg_11_53_inst : DFF_X1 port map( D => n7972, CK => clk, Q => 
                           n18462, QN => n2107);
   registers_reg_11_52_inst : DFF_X1 port map( D => n7971, CK => clk, Q => 
                           n18461, QN => n2108);
   registers_reg_11_51_inst : DFF_X1 port map( D => n7970, CK => clk, Q => 
                           n18460, QN => n2109);
   registers_reg_11_50_inst : DFF_X1 port map( D => n7969, CK => clk, Q => 
                           n18459, QN => n2110);
   registers_reg_11_49_inst : DFF_X1 port map( D => n7968, CK => clk, Q => 
                           n18458, QN => n2111);
   registers_reg_11_48_inst : DFF_X1 port map( D => n7967, CK => clk, Q => 
                           n18457, QN => n2112);
   registers_reg_11_47_inst : DFF_X1 port map( D => n7966, CK => clk, Q => 
                           n18456, QN => n2113);
   registers_reg_11_46_inst : DFF_X1 port map( D => n7965, CK => clk, Q => 
                           n18455, QN => n2114);
   registers_reg_11_45_inst : DFF_X1 port map( D => n7964, CK => clk, Q => 
                           n18454, QN => n2115);
   registers_reg_11_44_inst : DFF_X1 port map( D => n7963, CK => clk, Q => 
                           n18453, QN => n2116);
   registers_reg_11_43_inst : DFF_X1 port map( D => n7962, CK => clk, Q => 
                           n18452, QN => n2117);
   registers_reg_11_42_inst : DFF_X1 port map( D => n7961, CK => clk, Q => 
                           n18451, QN => n2118);
   registers_reg_11_41_inst : DFF_X1 port map( D => n7960, CK => clk, Q => 
                           n18450, QN => n2119);
   registers_reg_11_40_inst : DFF_X1 port map( D => n7959, CK => clk, Q => 
                           n18449, QN => n2120);
   registers_reg_11_39_inst : DFF_X1 port map( D => n7958, CK => clk, Q => 
                           n18448, QN => n2121);
   registers_reg_11_38_inst : DFF_X1 port map( D => n7957, CK => clk, Q => 
                           n18447, QN => n2122);
   registers_reg_11_37_inst : DFF_X1 port map( D => n7956, CK => clk, Q => 
                           n18446, QN => n2123);
   registers_reg_11_36_inst : DFF_X1 port map( D => n7955, CK => clk, Q => 
                           n18445, QN => n2124);
   registers_reg_11_35_inst : DFF_X1 port map( D => n7954, CK => clk, Q => 
                           n18444, QN => n2125);
   registers_reg_11_34_inst : DFF_X1 port map( D => n7953, CK => clk, Q => 
                           n18443, QN => n2126);
   registers_reg_11_33_inst : DFF_X1 port map( D => n7952, CK => clk, Q => 
                           n18442, QN => n2127);
   registers_reg_11_32_inst : DFF_X1 port map( D => n7951, CK => clk, Q => 
                           n18441, QN => n2128);
   registers_reg_11_31_inst : DFF_X1 port map( D => n7950, CK => clk, Q => 
                           n18440, QN => n2129);
   registers_reg_11_30_inst : DFF_X1 port map( D => n7949, CK => clk, Q => 
                           n18439, QN => n2130);
   registers_reg_11_29_inst : DFF_X1 port map( D => n7948, CK => clk, Q => 
                           n18438, QN => n2131);
   registers_reg_11_28_inst : DFF_X1 port map( D => n7947, CK => clk, Q => 
                           n18437, QN => n2132);
   registers_reg_11_27_inst : DFF_X1 port map( D => n7946, CK => clk, Q => 
                           n18436, QN => n2133);
   registers_reg_11_26_inst : DFF_X1 port map( D => n7945, CK => clk, Q => 
                           n18435, QN => n2134);
   registers_reg_11_25_inst : DFF_X1 port map( D => n7944, CK => clk, Q => 
                           n18434, QN => n2135);
   registers_reg_11_24_inst : DFF_X1 port map( D => n7943, CK => clk, Q => 
                           n18433, QN => n2136);
   registers_reg_11_23_inst : DFF_X1 port map( D => n7942, CK => clk, Q => 
                           n18432, QN => n2137);
   registers_reg_11_22_inst : DFF_X1 port map( D => n7941, CK => clk, Q => 
                           n18431, QN => n2138);
   registers_reg_11_21_inst : DFF_X1 port map( D => n7940, CK => clk, Q => 
                           n18430, QN => n2139);
   registers_reg_11_20_inst : DFF_X1 port map( D => n7939, CK => clk, Q => 
                           n18429, QN => n2140);
   registers_reg_11_19_inst : DFF_X1 port map( D => n7938, CK => clk, Q => 
                           n18428, QN => n2141);
   registers_reg_11_18_inst : DFF_X1 port map( D => n7937, CK => clk, Q => 
                           n18427, QN => n2142);
   registers_reg_11_17_inst : DFF_X1 port map( D => n7936, CK => clk, Q => 
                           n18426, QN => n2143);
   registers_reg_11_16_inst : DFF_X1 port map( D => n7935, CK => clk, Q => 
                           n18425, QN => n2144);
   registers_reg_11_15_inst : DFF_X1 port map( D => n7934, CK => clk, Q => 
                           n18424, QN => n2147);
   registers_reg_11_14_inst : DFF_X1 port map( D => n7933, CK => clk, Q => 
                           n18423, QN => n2150);
   registers_reg_11_13_inst : DFF_X1 port map( D => n7932, CK => clk, Q => 
                           n18422, QN => n2153);
   registers_reg_11_12_inst : DFF_X1 port map( D => n7931, CK => clk, Q => 
                           n18421, QN => n2156);
   registers_reg_11_11_inst : DFF_X1 port map( D => n7930, CK => clk, Q => 
                           n18420, QN => n2159);
   registers_reg_11_10_inst : DFF_X1 port map( D => n7929, CK => clk, Q => 
                           n18419, QN => n2162);
   registers_reg_11_9_inst : DFF_X1 port map( D => n7928, CK => clk, Q => 
                           n18418, QN => n2165);
   registers_reg_11_8_inst : DFF_X1 port map( D => n7927, CK => clk, Q => 
                           n18417, QN => n2168);
   registers_reg_11_7_inst : DFF_X1 port map( D => n7926, CK => clk, Q => 
                           n18416, QN => n2171);
   registers_reg_11_6_inst : DFF_X1 port map( D => n7925, CK => clk, Q => 
                           n18415, QN => n2174);
   registers_reg_11_5_inst : DFF_X1 port map( D => n7924, CK => clk, Q => 
                           n18414, QN => n2177);
   registers_reg_11_4_inst : DFF_X1 port map( D => n7923, CK => clk, Q => 
                           n18413, QN => n2180);
   registers_reg_4_63_inst : DFF_X1 port map( D => n7534, CK => clk, Q => 
                           registers_4_63_port, QN => n2261);
   registers_reg_4_62_inst : DFF_X1 port map( D => n7533, CK => clk, Q => 
                           registers_4_62_port, QN => n2264);
   registers_reg_4_61_inst : DFF_X1 port map( D => n7532, CK => clk, Q => 
                           registers_4_61_port, QN => n2267);
   registers_reg_4_60_inst : DFF_X1 port map( D => n7531, CK => clk, Q => 
                           registers_4_60_port, QN => n2270);
   registers_reg_4_59_inst : DFF_X1 port map( D => n7530, CK => clk, Q => 
                           registers_4_59_port, QN => n2273);
   registers_reg_4_58_inst : DFF_X1 port map( D => n7529, CK => clk, Q => 
                           registers_4_58_port, QN => n2276);
   registers_reg_4_57_inst : DFF_X1 port map( D => n7528, CK => clk, Q => 
                           registers_4_57_port, QN => n2279);
   registers_reg_4_56_inst : DFF_X1 port map( D => n7527, CK => clk, Q => 
                           registers_4_56_port, QN => n2282);
   registers_reg_4_55_inst : DFF_X1 port map( D => n7526, CK => clk, Q => 
                           registers_4_55_port, QN => n2285);
   registers_reg_4_54_inst : DFF_X1 port map( D => n7525, CK => clk, Q => 
                           registers_4_54_port, QN => n2288);
   registers_reg_4_53_inst : DFF_X1 port map( D => n7524, CK => clk, Q => 
                           registers_4_53_port, QN => n2291);
   registers_reg_4_52_inst : DFF_X1 port map( D => n7523, CK => clk, Q => 
                           registers_4_52_port, QN => n2294);
   registers_reg_4_51_inst : DFF_X1 port map( D => n7522, CK => clk, Q => 
                           registers_4_51_port, QN => n2297);
   registers_reg_4_50_inst : DFF_X1 port map( D => n7521, CK => clk, Q => 
                           registers_4_50_port, QN => n2300);
   registers_reg_4_49_inst : DFF_X1 port map( D => n7520, CK => clk, Q => 
                           registers_4_49_port, QN => n2303);
   registers_reg_4_48_inst : DFF_X1 port map( D => n7519, CK => clk, Q => 
                           registers_4_48_port, QN => n2306);
   registers_reg_4_47_inst : DFF_X1 port map( D => n7518, CK => clk, Q => 
                           registers_4_47_port, QN => n2309);
   registers_reg_4_46_inst : DFF_X1 port map( D => n7517, CK => clk, Q => 
                           registers_4_46_port, QN => n2312);
   registers_reg_4_45_inst : DFF_X1 port map( D => n7516, CK => clk, Q => 
                           registers_4_45_port, QN => n2315);
   registers_reg_4_44_inst : DFF_X1 port map( D => n7515, CK => clk, Q => 
                           registers_4_44_port, QN => n2318);
   registers_reg_4_43_inst : DFF_X1 port map( D => n7514, CK => clk, Q => 
                           registers_4_43_port, QN => n2321);
   registers_reg_4_42_inst : DFF_X1 port map( D => n7513, CK => clk, Q => 
                           registers_4_42_port, QN => n2324);
   registers_reg_4_41_inst : DFF_X1 port map( D => n7512, CK => clk, Q => 
                           registers_4_41_port, QN => n2327);
   registers_reg_4_40_inst : DFF_X1 port map( D => n7511, CK => clk, Q => 
                           registers_4_40_port, QN => n2330);
   registers_reg_4_39_inst : DFF_X1 port map( D => n7510, CK => clk, Q => 
                           registers_4_39_port, QN => n2333);
   registers_reg_4_38_inst : DFF_X1 port map( D => n7509, CK => clk, Q => 
                           registers_4_38_port, QN => n2336);
   registers_reg_4_37_inst : DFF_X1 port map( D => n7508, CK => clk, Q => 
                           registers_4_37_port, QN => n2337);
   registers_reg_4_36_inst : DFF_X1 port map( D => n7507, CK => clk, Q => 
                           registers_4_36_port, QN => n2338);
   registers_reg_4_35_inst : DFF_X1 port map( D => n7506, CK => clk, Q => 
                           registers_4_35_port, QN => n2339);
   registers_reg_4_34_inst : DFF_X1 port map( D => n7505, CK => clk, Q => 
                           registers_4_34_port, QN => n2340);
   registers_reg_4_33_inst : DFF_X1 port map( D => n7504, CK => clk, Q => 
                           registers_4_33_port, QN => n2341);
   registers_reg_4_32_inst : DFF_X1 port map( D => n7503, CK => clk, Q => 
                           registers_4_32_port, QN => n2342);
   registers_reg_4_31_inst : DFF_X1 port map( D => n7502, CK => clk, Q => 
                           registers_4_31_port, QN => n2343);
   registers_reg_4_30_inst : DFF_X1 port map( D => n7501, CK => clk, Q => 
                           registers_4_30_port, QN => n2344);
   registers_reg_4_29_inst : DFF_X1 port map( D => n7500, CK => clk, Q => 
                           registers_4_29_port, QN => n2345);
   registers_reg_4_28_inst : DFF_X1 port map( D => n7499, CK => clk, Q => 
                           registers_4_28_port, QN => n2346);
   registers_reg_4_27_inst : DFF_X1 port map( D => n7498, CK => clk, Q => 
                           registers_4_27_port, QN => n2347);
   registers_reg_4_26_inst : DFF_X1 port map( D => n7497, CK => clk, Q => 
                           registers_4_26_port, QN => n2348);
   registers_reg_4_25_inst : DFF_X1 port map( D => n7496, CK => clk, Q => 
                           registers_4_25_port, QN => n2349);
   registers_reg_4_24_inst : DFF_X1 port map( D => n7495, CK => clk, Q => 
                           registers_4_24_port, QN => n2350);
   registers_reg_4_23_inst : DFF_X1 port map( D => n7494, CK => clk, Q => 
                           registers_4_23_port, QN => n2351);
   registers_reg_4_22_inst : DFF_X1 port map( D => n7493, CK => clk, Q => 
                           registers_4_22_port, QN => n2352);
   registers_reg_4_21_inst : DFF_X1 port map( D => n7492, CK => clk, Q => 
                           registers_4_21_port, QN => n2353);
   registers_reg_4_20_inst : DFF_X1 port map( D => n7491, CK => clk, Q => 
                           registers_4_20_port, QN => n2354);
   registers_reg_4_19_inst : DFF_X1 port map( D => n7490, CK => clk, Q => 
                           registers_4_19_port, QN => n2355);
   registers_reg_4_18_inst : DFF_X1 port map( D => n7489, CK => clk, Q => 
                           registers_4_18_port, QN => n2356);
   registers_reg_4_17_inst : DFF_X1 port map( D => n7488, CK => clk, Q => 
                           registers_4_17_port, QN => n2357);
   registers_reg_4_16_inst : DFF_X1 port map( D => n7487, CK => clk, Q => 
                           registers_4_16_port, QN => n2358);
   registers_reg_4_15_inst : DFF_X1 port map( D => n7486, CK => clk, Q => 
                           registers_4_15_port, QN => n2359);
   registers_reg_4_14_inst : DFF_X1 port map( D => n7485, CK => clk, Q => 
                           registers_4_14_port, QN => n2360);
   registers_reg_4_13_inst : DFF_X1 port map( D => n7484, CK => clk, Q => 
                           registers_4_13_port, QN => n2361);
   registers_reg_4_12_inst : DFF_X1 port map( D => n7483, CK => clk, Q => 
                           registers_4_12_port, QN => n2362);
   registers_reg_4_11_inst : DFF_X1 port map( D => n7482, CK => clk, Q => 
                           registers_4_11_port, QN => n2363);
   registers_reg_4_10_inst : DFF_X1 port map( D => n7481, CK => clk, Q => 
                           registers_4_10_port, QN => n2364);
   registers_reg_4_9_inst : DFF_X1 port map( D => n7480, CK => clk, Q => 
                           registers_4_9_port, QN => n2365);
   registers_reg_4_8_inst : DFF_X1 port map( D => n7479, CK => clk, Q => 
                           registers_4_8_port, QN => n2366);
   registers_reg_4_7_inst : DFF_X1 port map( D => n7478, CK => clk, Q => 
                           registers_4_7_port, QN => n2367);
   registers_reg_4_6_inst : DFF_X1 port map( D => n7477, CK => clk, Q => 
                           registers_4_6_port, QN => n2368);
   registers_reg_4_5_inst : DFF_X1 port map( D => n7476, CK => clk, Q => 
                           registers_4_5_port, QN => n2369);
   registers_reg_4_4_inst : DFF_X1 port map( D => n7475, CK => clk, Q => 
                           registers_4_4_port, QN => n2370);
   registers_reg_22_63_inst : DFF_X1 port map( D => n8686, CK => clk, Q => 
                           n18412, QN => n1730);
   registers_reg_22_62_inst : DFF_X1 port map( D => n8685, CK => clk, Q => 
                           n18411, QN => n1731);
   registers_reg_22_61_inst : DFF_X1 port map( D => n8684, CK => clk, Q => 
                           n18410, QN => n1732);
   registers_reg_22_60_inst : DFF_X1 port map( D => n8683, CK => clk, Q => 
                           n18409, QN => n1733);
   registers_reg_22_59_inst : DFF_X1 port map( D => n8682, CK => clk, Q => 
                           n18408, QN => n1734);
   registers_reg_22_58_inst : DFF_X1 port map( D => n8681, CK => clk, Q => 
                           n18407, QN => n1735);
   registers_reg_22_57_inst : DFF_X1 port map( D => n8680, CK => clk, Q => 
                           n18406, QN => n1736);
   registers_reg_22_56_inst : DFF_X1 port map( D => n8679, CK => clk, Q => 
                           n18405, QN => n1737);
   registers_reg_22_55_inst : DFF_X1 port map( D => n8678, CK => clk, Q => 
                           n18404, QN => n1738);
   registers_reg_22_54_inst : DFF_X1 port map( D => n8677, CK => clk, Q => 
                           n18403, QN => n1739);
   registers_reg_22_53_inst : DFF_X1 port map( D => n8676, CK => clk, Q => 
                           n18402, QN => n1740);
   registers_reg_22_52_inst : DFF_X1 port map( D => n8675, CK => clk, Q => 
                           n18401, QN => n1741);
   registers_reg_22_51_inst : DFF_X1 port map( D => n8674, CK => clk, Q => 
                           n18400, QN => n1742);
   registers_reg_22_50_inst : DFF_X1 port map( D => n8673, CK => clk, Q => 
                           n18399, QN => n1743);
   registers_reg_22_49_inst : DFF_X1 port map( D => n8672, CK => clk, Q => 
                           n18398, QN => n1744);
   registers_reg_22_48_inst : DFF_X1 port map( D => n8671, CK => clk, Q => 
                           n18397, QN => n1745);
   registers_reg_22_47_inst : DFF_X1 port map( D => n8670, CK => clk, Q => 
                           n18396, QN => n1749);
   registers_reg_22_46_inst : DFF_X1 port map( D => n8669, CK => clk, Q => 
                           n18395, QN => n1750);
   registers_reg_22_45_inst : DFF_X1 port map( D => n8668, CK => clk, Q => 
                           n18394, QN => n1751);
   registers_reg_22_44_inst : DFF_X1 port map( D => n8667, CK => clk, Q => 
                           n18393, QN => n1752);
   registers_reg_22_43_inst : DFF_X1 port map( D => n8666, CK => clk, Q => 
                           n18392, QN => n1753);
   registers_reg_22_42_inst : DFF_X1 port map( D => n8665, CK => clk, Q => 
                           n18391, QN => n1754);
   registers_reg_22_41_inst : DFF_X1 port map( D => n8664, CK => clk, Q => 
                           n18390, QN => n1755);
   registers_reg_22_40_inst : DFF_X1 port map( D => n8663, CK => clk, Q => 
                           n18389, QN => n1756);
   registers_reg_22_39_inst : DFF_X1 port map( D => n8662, CK => clk, Q => 
                           n18388, QN => n1757);
   registers_reg_22_38_inst : DFF_X1 port map( D => n8661, CK => clk, Q => 
                           n18387, QN => n1758);
   registers_reg_22_37_inst : DFF_X1 port map( D => n8660, CK => clk, Q => 
                           n18386, QN => n1759);
   registers_reg_22_36_inst : DFF_X1 port map( D => n8659, CK => clk, Q => 
                           n18385, QN => n1760);
   registers_reg_22_35_inst : DFF_X1 port map( D => n8658, CK => clk, Q => 
                           n18384, QN => n1761);
   registers_reg_22_34_inst : DFF_X1 port map( D => n8657, CK => clk, Q => 
                           n18383, QN => n1762);
   registers_reg_22_33_inst : DFF_X1 port map( D => n8656, CK => clk, Q => 
                           n18382, QN => n1763);
   registers_reg_22_32_inst : DFF_X1 port map( D => n8655, CK => clk, Q => 
                           n18381, QN => n1764);
   registers_reg_22_31_inst : DFF_X1 port map( D => n8654, CK => clk, Q => 
                           n18380, QN => n1765);
   registers_reg_22_30_inst : DFF_X1 port map( D => n8653, CK => clk, Q => 
                           n18379, QN => n1766);
   registers_reg_22_29_inst : DFF_X1 port map( D => n8652, CK => clk, Q => 
                           n18378, QN => n1767);
   registers_reg_22_28_inst : DFF_X1 port map( D => n8651, CK => clk, Q => 
                           n18377, QN => n1768);
   registers_reg_22_27_inst : DFF_X1 port map( D => n8650, CK => clk, Q => 
                           n18376, QN => n1769);
   registers_reg_22_26_inst : DFF_X1 port map( D => n8649, CK => clk, Q => 
                           n18375, QN => n1770);
   registers_reg_22_25_inst : DFF_X1 port map( D => n8648, CK => clk, Q => 
                           n18374, QN => n1771);
   registers_reg_22_24_inst : DFF_X1 port map( D => n8647, CK => clk, Q => 
                           n18373, QN => n1772);
   registers_reg_22_23_inst : DFF_X1 port map( D => n8646, CK => clk, Q => 
                           n18372, QN => n1773);
   registers_reg_22_22_inst : DFF_X1 port map( D => n8645, CK => clk, Q => 
                           n18371, QN => n1774);
   registers_reg_22_21_inst : DFF_X1 port map( D => n8644, CK => clk, Q => 
                           n18370, QN => n1775);
   registers_reg_22_20_inst : DFF_X1 port map( D => n8643, CK => clk, Q => 
                           n18369, QN => n1776);
   registers_reg_22_19_inst : DFF_X1 port map( D => n8642, CK => clk, Q => 
                           n18368, QN => n1777);
   registers_reg_22_18_inst : DFF_X1 port map( D => n8641, CK => clk, Q => 
                           n18367, QN => n1778);
   registers_reg_22_17_inst : DFF_X1 port map( D => n8640, CK => clk, Q => 
                           n18366, QN => n1779);
   registers_reg_22_16_inst : DFF_X1 port map( D => n8639, CK => clk, Q => 
                           n18365, QN => n1780);
   registers_reg_22_15_inst : DFF_X1 port map( D => n8638, CK => clk, Q => 
                           n18364, QN => n1781);
   registers_reg_22_14_inst : DFF_X1 port map( D => n8637, CK => clk, Q => 
                           n18363, QN => n1782);
   registers_reg_22_13_inst : DFF_X1 port map( D => n8636, CK => clk, Q => 
                           n18362, QN => n1783);
   registers_reg_22_12_inst : DFF_X1 port map( D => n8635, CK => clk, Q => 
                           n18361, QN => n1784);
   registers_reg_22_11_inst : DFF_X1 port map( D => n8634, CK => clk, Q => 
                           n18360, QN => n1785);
   registers_reg_22_10_inst : DFF_X1 port map( D => n8633, CK => clk, Q => 
                           n18359, QN => n1786);
   registers_reg_22_9_inst : DFF_X1 port map( D => n8632, CK => clk, Q => 
                           n18358, QN => n1787);
   registers_reg_22_8_inst : DFF_X1 port map( D => n8631, CK => clk, Q => 
                           n18357, QN => n1788);
   registers_reg_22_7_inst : DFF_X1 port map( D => n8630, CK => clk, Q => 
                           n18356, QN => n1789);
   registers_reg_22_6_inst : DFF_X1 port map( D => n8629, CK => clk, Q => 
                           n18355, QN => n1790);
   registers_reg_22_5_inst : DFF_X1 port map( D => n8628, CK => clk, Q => 
                           n18354, QN => n1791);
   registers_reg_22_4_inst : DFF_X1 port map( D => n8627, CK => clk, Q => 
                           n18353, QN => n1792);
   out_to_mem_reg_47_inst : DFF_X1 port map( D => n7211, CK => clk, Q => 
                           out_to_mem_47_port, QN => n18352);
   out_to_mem_reg_46_inst : DFF_X1 port map( D => n7207, CK => clk, Q => 
                           out_to_mem_46_port, QN => n18351);
   out_to_mem_reg_45_inst : DFF_X1 port map( D => n7203, CK => clk, Q => 
                           out_to_mem_45_port, QN => n18350);
   out_to_mem_reg_44_inst : DFF_X1 port map( D => n7199, CK => clk, Q => 
                           out_to_mem_44_port, QN => n18349);
   out_to_mem_reg_43_inst : DFF_X1 port map( D => n7195, CK => clk, Q => 
                           out_to_mem_43_port, QN => n18348);
   out_to_mem_reg_42_inst : DFF_X1 port map( D => n7191, CK => clk, Q => 
                           out_to_mem_42_port, QN => n18347);
   out_to_mem_reg_41_inst : DFF_X1 port map( D => n7187, CK => clk, Q => 
                           out_to_mem_41_port, QN => n18346);
   out_to_mem_reg_40_inst : DFF_X1 port map( D => n7183, CK => clk, Q => 
                           out_to_mem_40_port, QN => n18345);
   out_to_mem_reg_39_inst : DFF_X1 port map( D => n7179, CK => clk, Q => 
                           out_to_mem_39_port, QN => n18344);
   out_to_mem_reg_38_inst : DFF_X1 port map( D => n7175, CK => clk, Q => 
                           out_to_mem_38_port, QN => n18343);
   out_to_mem_reg_37_inst : DFF_X1 port map( D => n7171, CK => clk, Q => 
                           out_to_mem_37_port, QN => n18342);
   out_to_mem_reg_36_inst : DFF_X1 port map( D => n7167, CK => clk, Q => 
                           out_to_mem_36_port, QN => n18341);
   registers_reg_21_63_inst : DFF_X1 port map( D => n8622, CK => clk, Q => 
                           n18340, QN => n1800);
   registers_reg_21_62_inst : DFF_X1 port map( D => n8621, CK => clk, Q => 
                           n18339, QN => n1801);
   registers_reg_21_61_inst : DFF_X1 port map( D => n8620, CK => clk, Q => 
                           n18338, QN => n1802);
   registers_reg_21_60_inst : DFF_X1 port map( D => n8619, CK => clk, Q => 
                           n18337, QN => n1803);
   registers_reg_21_59_inst : DFF_X1 port map( D => n8618, CK => clk, Q => 
                           n18336, QN => n1804);
   registers_reg_21_58_inst : DFF_X1 port map( D => n8617, CK => clk, Q => 
                           n18335, QN => n1805);
   registers_reg_21_57_inst : DFF_X1 port map( D => n8616, CK => clk, Q => 
                           n18334, QN => n1806);
   registers_reg_21_56_inst : DFF_X1 port map( D => n8615, CK => clk, Q => 
                           n18333, QN => n1807);
   registers_reg_21_55_inst : DFF_X1 port map( D => n8614, CK => clk, Q => 
                           n18332, QN => n1808);
   registers_reg_21_54_inst : DFF_X1 port map( D => n8613, CK => clk, Q => 
                           n18331, QN => n1809);
   registers_reg_21_53_inst : DFF_X1 port map( D => n8612, CK => clk, Q => 
                           n18330, QN => n1810);
   registers_reg_21_52_inst : DFF_X1 port map( D => n8611, CK => clk, Q => 
                           n18329, QN => n1811);
   registers_reg_21_51_inst : DFF_X1 port map( D => n8610, CK => clk, Q => 
                           n18328, QN => n1812);
   registers_reg_21_50_inst : DFF_X1 port map( D => n8609, CK => clk, Q => 
                           n18327, QN => n1813);
   registers_reg_21_49_inst : DFF_X1 port map( D => n8608, CK => clk, Q => 
                           n18326, QN => n1814);
   registers_reg_21_48_inst : DFF_X1 port map( D => n8607, CK => clk, Q => 
                           n18325, QN => n1815);
   registers_reg_21_47_inst : DFF_X1 port map( D => n8606, CK => clk, Q => 
                           n18324, QN => n1816);
   registers_reg_21_46_inst : DFF_X1 port map( D => n8605, CK => clk, Q => 
                           n18323, QN => n1817);
   registers_reg_21_45_inst : DFF_X1 port map( D => n8604, CK => clk, Q => 
                           n18322, QN => n1818);
   registers_reg_21_44_inst : DFF_X1 port map( D => n8603, CK => clk, Q => 
                           n18321, QN => n1819);
   registers_reg_21_43_inst : DFF_X1 port map( D => n8602, CK => clk, Q => 
                           n18320, QN => n1820);
   registers_reg_21_42_inst : DFF_X1 port map( D => n8601, CK => clk, Q => 
                           n18319, QN => n1821);
   registers_reg_21_41_inst : DFF_X1 port map( D => n8600, CK => clk, Q => 
                           n18318, QN => n1822);
   registers_reg_21_40_inst : DFF_X1 port map( D => n8599, CK => clk, Q => 
                           n18317, QN => n1823);
   registers_reg_21_39_inst : DFF_X1 port map( D => n8598, CK => clk, Q => 
                           n18316, QN => n1824);
   registers_reg_21_38_inst : DFF_X1 port map( D => n8597, CK => clk, Q => 
                           n18315, QN => n1825);
   registers_reg_21_37_inst : DFF_X1 port map( D => n8596, CK => clk, Q => 
                           n18314, QN => n1826);
   registers_reg_21_36_inst : DFF_X1 port map( D => n8595, CK => clk, Q => 
                           n18313, QN => n1827);
   registers_reg_21_35_inst : DFF_X1 port map( D => n8594, CK => clk, Q => 
                           n18312, QN => n1828);
   registers_reg_21_34_inst : DFF_X1 port map( D => n8593, CK => clk, Q => 
                           n18311, QN => n1829);
   registers_reg_21_33_inst : DFF_X1 port map( D => n8592, CK => clk, Q => 
                           n18310, QN => n1830);
   registers_reg_21_32_inst : DFF_X1 port map( D => n8591, CK => clk, Q => 
                           n18309, QN => n1831);
   registers_reg_21_31_inst : DFF_X1 port map( D => n8590, CK => clk, Q => 
                           n18308, QN => n1832);
   registers_reg_21_30_inst : DFF_X1 port map( D => n8589, CK => clk, Q => 
                           n18307, QN => n1833);
   registers_reg_21_29_inst : DFF_X1 port map( D => n8588, CK => clk, Q => 
                           n18306, QN => n1834);
   registers_reg_21_28_inst : DFF_X1 port map( D => n8587, CK => clk, Q => 
                           n18305, QN => n1835);
   registers_reg_21_27_inst : DFF_X1 port map( D => n8586, CK => clk, Q => 
                           n18304, QN => n1836);
   registers_reg_21_26_inst : DFF_X1 port map( D => n8585, CK => clk, Q => 
                           n18303, QN => n1837);
   registers_reg_21_25_inst : DFF_X1 port map( D => n8584, CK => clk, Q => 
                           n18302, QN => n1838);
   registers_reg_21_24_inst : DFF_X1 port map( D => n8583, CK => clk, Q => 
                           n18301, QN => n1839);
   registers_reg_21_23_inst : DFF_X1 port map( D => n8582, CK => clk, Q => 
                           n18300, QN => n1840);
   registers_reg_21_22_inst : DFF_X1 port map( D => n8581, CK => clk, Q => 
                           n18299, QN => n1841);
   registers_reg_21_21_inst : DFF_X1 port map( D => n8580, CK => clk, Q => 
                           n18298, QN => n1842);
   registers_reg_21_20_inst : DFF_X1 port map( D => n8579, CK => clk, Q => 
                           n18297, QN => n1843);
   registers_reg_21_19_inst : DFF_X1 port map( D => n8578, CK => clk, Q => 
                           n18296, QN => n1844);
   registers_reg_21_18_inst : DFF_X1 port map( D => n8577, CK => clk, Q => 
                           n18295, QN => n1845);
   registers_reg_21_17_inst : DFF_X1 port map( D => n8576, CK => clk, Q => 
                           n18294, QN => n1846);
   registers_reg_21_16_inst : DFF_X1 port map( D => n8575, CK => clk, Q => 
                           n18293, QN => n1847);
   registers_reg_21_15_inst : DFF_X1 port map( D => n8574, CK => clk, Q => 
                           n18292, QN => n1848);
   registers_reg_21_14_inst : DFF_X1 port map( D => n8573, CK => clk, Q => 
                           n18291, QN => n1849);
   registers_reg_21_13_inst : DFF_X1 port map( D => n8572, CK => clk, Q => 
                           n18290, QN => n1850);
   registers_reg_21_12_inst : DFF_X1 port map( D => n8571, CK => clk, Q => 
                           n18289, QN => n1851);
   registers_reg_21_11_inst : DFF_X1 port map( D => n8570, CK => clk, Q => 
                           n18288, QN => n1852);
   registers_reg_21_10_inst : DFF_X1 port map( D => n8569, CK => clk, Q => 
                           n18287, QN => n1853);
   registers_reg_21_9_inst : DFF_X1 port map( D => n8568, CK => clk, Q => 
                           n18286, QN => n1854);
   registers_reg_21_8_inst : DFF_X1 port map( D => n8567, CK => clk, Q => 
                           n18285, QN => n1855);
   registers_reg_21_7_inst : DFF_X1 port map( D => n8566, CK => clk, Q => 
                           n18284, QN => n1856);
   registers_reg_21_6_inst : DFF_X1 port map( D => n8565, CK => clk, Q => 
                           n18283, QN => n1857);
   registers_reg_21_5_inst : DFF_X1 port map( D => n8564, CK => clk, Q => 
                           n18282, QN => n1858);
   registers_reg_21_4_inst : DFF_X1 port map( D => n8563, CK => clk, Q => 
                           n18281, QN => n1859);
   out_to_mem_reg_59_inst : DFF_X1 port map( D => n7259, CK => clk, Q => 
                           out_to_mem_59_port, QN => n18280);
   out_to_mem_reg_58_inst : DFF_X1 port map( D => n7255, CK => clk, Q => 
                           out_to_mem_58_port, QN => n18279);
   out_to_mem_reg_57_inst : DFF_X1 port map( D => n7251, CK => clk, Q => 
                           out_to_mem_57_port, QN => n18278);
   out_to_mem_reg_56_inst : DFF_X1 port map( D => n7247, CK => clk, Q => 
                           out_to_mem_56_port, QN => n18277);
   out_to_mem_reg_55_inst : DFF_X1 port map( D => n7243, CK => clk, Q => 
                           out_to_mem_55_port, QN => n18276);
   out_to_mem_reg_54_inst : DFF_X1 port map( D => n7239, CK => clk, Q => 
                           out_to_mem_54_port, QN => n18275);
   out_to_mem_reg_53_inst : DFF_X1 port map( D => n7235, CK => clk, Q => 
                           out_to_mem_53_port, QN => n18274);
   out_to_mem_reg_52_inst : DFF_X1 port map( D => n7231, CK => clk, Q => 
                           out_to_mem_52_port, QN => n18273);
   out_to_mem_reg_51_inst : DFF_X1 port map( D => n7227, CK => clk, Q => 
                           out_to_mem_51_port, QN => n18272);
   out_to_mem_reg_50_inst : DFF_X1 port map( D => n7223, CK => clk, Q => 
                           out_to_mem_50_port, QN => n18271);
   out_to_mem_reg_49_inst : DFF_X1 port map( D => n7219, CK => clk, Q => 
                           out_to_mem_49_port, QN => n18270);
   out_to_mem_reg_48_inst : DFF_X1 port map( D => n7215, CK => clk, Q => 
                           out_to_mem_48_port, QN => n18269);
   out_to_mem_reg_35_inst : DFF_X1 port map( D => n7163, CK => clk, Q => 
                           out_to_mem_35_port, QN => n18268);
   out_to_mem_reg_34_inst : DFF_X1 port map( D => n7159, CK => clk, Q => 
                           out_to_mem_34_port, QN => n18267);
   out_to_mem_reg_33_inst : DFF_X1 port map( D => n7155, CK => clk, Q => 
                           out_to_mem_33_port, QN => n18266);
   out_to_mem_reg_32_inst : DFF_X1 port map( D => n7151, CK => clk, Q => 
                           out_to_mem_32_port, QN => n18265);
   out_to_mem_reg_31_inst : DFF_X1 port map( D => n7147, CK => clk, Q => 
                           out_to_mem_31_port, QN => n18264);
   out_to_mem_reg_30_inst : DFF_X1 port map( D => n7143, CK => clk, Q => 
                           out_to_mem_30_port, QN => n18263);
   out_to_mem_reg_29_inst : DFF_X1 port map( D => n7139, CK => clk, Q => 
                           out_to_mem_29_port, QN => n18262);
   out_to_mem_reg_28_inst : DFF_X1 port map( D => n7135, CK => clk, Q => 
                           out_to_mem_28_port, QN => n18261);
   out_to_mem_reg_27_inst : DFF_X1 port map( D => n7131, CK => clk, Q => 
                           out_to_mem_27_port, QN => n18260);
   out_to_mem_reg_26_inst : DFF_X1 port map( D => n7127, CK => clk, Q => 
                           out_to_mem_26_port, QN => n18259);
   out_to_mem_reg_25_inst : DFF_X1 port map( D => n7123, CK => clk, Q => 
                           out_to_mem_25_port, QN => n18258);
   out_to_mem_reg_24_inst : DFF_X1 port map( D => n7119, CK => clk, Q => 
                           out_to_mem_24_port, QN => n18257);
   out_to_mem_reg_23_inst : DFF_X1 port map( D => n7115, CK => clk, Q => 
                           out_to_mem_23_port, QN => n18256);
   out_to_mem_reg_22_inst : DFF_X1 port map( D => n7111, CK => clk, Q => 
                           out_to_mem_22_port, QN => n18255);
   out_to_mem_reg_21_inst : DFF_X1 port map( D => n7107, CK => clk, Q => 
                           out_to_mem_21_port, QN => n18254);
   out_to_mem_reg_20_inst : DFF_X1 port map( D => n7103, CK => clk, Q => 
                           out_to_mem_20_port, QN => n18253);
   out_to_mem_reg_19_inst : DFF_X1 port map( D => n7099, CK => clk, Q => 
                           out_to_mem_19_port, QN => n18252);
   out_to_mem_reg_18_inst : DFF_X1 port map( D => n7095, CK => clk, Q => 
                           out_to_mem_18_port, QN => n18251);
   out_to_mem_reg_17_inst : DFF_X1 port map( D => n7091, CK => clk, Q => 
                           out_to_mem_17_port, QN => n18250);
   out_to_mem_reg_16_inst : DFF_X1 port map( D => n7087, CK => clk, Q => 
                           out_to_mem_16_port, QN => n18249);
   out_to_mem_reg_15_inst : DFF_X1 port map( D => n7083, CK => clk, Q => 
                           out_to_mem_15_port, QN => n18248);
   out_to_mem_reg_14_inst : DFF_X1 port map( D => n7079, CK => clk, Q => 
                           out_to_mem_14_port, QN => n18247);
   out_to_mem_reg_13_inst : DFF_X1 port map( D => n7075, CK => clk, Q => 
                           out_to_mem_13_port, QN => n18246);
   out_to_mem_reg_12_inst : DFF_X1 port map( D => n7071, CK => clk, Q => 
                           out_to_mem_12_port, QN => n18245);
   out_to_mem_reg_11_inst : DFF_X1 port map( D => n7067, CK => clk, Q => 
                           out_to_mem_11_port, QN => n18244);
   out_to_mem_reg_10_inst : DFF_X1 port map( D => n7063, CK => clk, Q => 
                           out_to_mem_10_port, QN => n18243);
   out_to_mem_reg_9_inst : DFF_X1 port map( D => n7059, CK => clk, Q => 
                           out_to_mem_9_port, QN => n18242);
   out_to_mem_reg_8_inst : DFF_X1 port map( D => n7055, CK => clk, Q => 
                           out_to_mem_8_port, QN => n18241);
   out_to_mem_reg_7_inst : DFF_X1 port map( D => n7051, CK => clk, Q => 
                           out_to_mem_7_port, QN => n18240);
   out_to_mem_reg_6_inst : DFF_X1 port map( D => n7047, CK => clk, Q => 
                           out_to_mem_6_port, QN => n18239);
   out_to_mem_reg_5_inst : DFF_X1 port map( D => n7043, CK => clk, Q => 
                           out_to_mem_5_port, QN => n18238);
   out_to_mem_reg_4_inst : DFF_X1 port map( D => n7039, CK => clk, Q => 
                           out_to_mem_4_port, QN => n18237);
   out_to_mem_reg_3_inst : DFF_X1 port map( D => n7035, CK => clk, Q => 
                           out_to_mem_3_port, QN => n18236);
   U3 : XOR2_X1 port map( A => n11725, B => n11726, Z => n1946);
   U4 : AOI21_X1 port map( B1 => add_wr(3), B2 => n11756, A => add_wr(4), ZN =>
                           n11751);
   U5 : AOI21_X1 port map( B1 => add_rd1(3), B2 => n11758, A => add_rd1(4), ZN 
                           => n11752);
   U9 : NAND3_X1 port map( A1 => count3(0), A2 => n1946, A3 => n1943, ZN => 
                           n2086);
   U10 : OAI21_X1 port map( B1 => U3_U2_Z_0, B2 => n11749, A => 
                           sub_86_carry_4_port, ZN => n11656);
   U11 : AOI21_X1 port map( B1 => n11752, B2 => sub_86_carry_4_port, A => 
                           n11749, ZN => n11654);
   U12 : INV_X1 port map( A => n11693, ZN => n3160);
   U13 : OAI22_X1 port map( A1 => n2375, A2 => n11709, B1 => n11695, B2 => 
                           n11710, ZN => n3166);
   U14 : BUF_X1 port map( A => n19489, Z => n19511);
   U15 : BUF_X1 port map( A => n19825, Z => n19847);
   U16 : BUF_X1 port map( A => n19713, Z => n19735);
   U17 : BUF_X1 port map( A => n19601, Z => n19623);
   U18 : BUF_X1 port map( A => n20049, Z => n20071);
   U19 : BUF_X1 port map( A => n20105, Z => n20127);
   U20 : BUF_X1 port map( A => n19657, Z => n19679);
   U21 : BUF_X1 port map( A => n20273, Z => n20295);
   U22 : BUF_X1 port map( A => n19937, Z => n19959);
   U23 : BUF_X1 port map( A => n20161, Z => n20183);
   U24 : BUF_X1 port map( A => n19881, Z => n19903);
   U25 : BUF_X1 port map( A => n19769, Z => n19791);
   U26 : BUF_X1 port map( A => n19545, Z => n19567);
   U27 : BUF_X1 port map( A => n20329, Z => n20351);
   U28 : BUF_X1 port map( A => n19993, Z => n20015);
   U29 : BUF_X1 port map( A => n20217, Z => n20239);
   U30 : BUF_X1 port map( A => n19573, Z => n19595);
   U31 : BUF_X1 port map( A => n19797, Z => n19819);
   U32 : BUF_X1 port map( A => n19685, Z => n19707);
   U33 : BUF_X1 port map( A => n19909, Z => n19931);
   U34 : BUF_X1 port map( A => n20133, Z => n20155);
   U35 : BUF_X1 port map( A => n20077, Z => n20099);
   U36 : BUF_X1 port map( A => n19629, Z => n19651);
   U37 : BUF_X1 port map( A => n20301, Z => n20323);
   U38 : BUF_X1 port map( A => n19965, Z => n19987);
   U39 : BUF_X1 port map( A => n20189, Z => n20211);
   U40 : BUF_X1 port map( A => n19517, Z => n19539);
   U41 : BUF_X1 port map( A => n19741, Z => n19763);
   U42 : BUF_X1 port map( A => n19853, Z => n19875);
   U43 : BUF_X1 port map( A => n20021, Z => n20043);
   U44 : BUF_X1 port map( A => n20549, Z => n20571);
   U45 : BUF_X1 port map( A => n20245, Z => n20267);
   U46 : INV_X1 port map( A => n19847, ZN => n19830);
   U47 : INV_X1 port map( A => n19847, ZN => n19829);
   U48 : INV_X1 port map( A => n19847, ZN => n19828);
   U49 : INV_X1 port map( A => n19735, ZN => n19718);
   U50 : INV_X1 port map( A => n19735, ZN => n19717);
   U51 : INV_X1 port map( A => n19735, ZN => n19716);
   U52 : INV_X1 port map( A => n19623, ZN => n19606);
   U53 : INV_X1 port map( A => n19623, ZN => n19605);
   U54 : INV_X1 port map( A => n19623, ZN => n19604);
   U55 : INV_X1 port map( A => n20071, ZN => n20054);
   U56 : INV_X1 port map( A => n20071, ZN => n20053);
   U57 : INV_X1 port map( A => n20071, ZN => n20052);
   U58 : INV_X1 port map( A => n20127, ZN => n20110);
   U59 : INV_X1 port map( A => n20127, ZN => n20109);
   U60 : INV_X1 port map( A => n20127, ZN => n20108);
   U61 : INV_X1 port map( A => n19679, ZN => n19662);
   U62 : INV_X1 port map( A => n19679, ZN => n19661);
   U63 : INV_X1 port map( A => n19679, ZN => n19660);
   U64 : INV_X1 port map( A => n20295, ZN => n20278);
   U65 : INV_X1 port map( A => n20295, ZN => n20277);
   U66 : INV_X1 port map( A => n20295, ZN => n20276);
   U67 : INV_X1 port map( A => n19959, ZN => n19942);
   U68 : INV_X1 port map( A => n19959, ZN => n19941);
   U69 : INV_X1 port map( A => n19959, ZN => n19940);
   U70 : INV_X1 port map( A => n20183, ZN => n20166);
   U71 : INV_X1 port map( A => n20183, ZN => n20165);
   U72 : INV_X1 port map( A => n20183, ZN => n20164);
   U73 : INV_X1 port map( A => n19903, ZN => n19886);
   U74 : INV_X1 port map( A => n19903, ZN => n19885);
   U75 : INV_X1 port map( A => n19903, ZN => n19884);
   U76 : INV_X1 port map( A => n19791, ZN => n19774);
   U77 : INV_X1 port map( A => n19791, ZN => n19773);
   U78 : INV_X1 port map( A => n19791, ZN => n19772);
   U79 : INV_X1 port map( A => n19567, ZN => n19550);
   U80 : INV_X1 port map( A => n19567, ZN => n19549);
   U81 : INV_X1 port map( A => n19567, ZN => n19548);
   U82 : INV_X1 port map( A => n20351, ZN => n20334);
   U83 : INV_X1 port map( A => n20351, ZN => n20333);
   U84 : INV_X1 port map( A => n20351, ZN => n20332);
   U85 : INV_X1 port map( A => n20015, ZN => n19998);
   U86 : INV_X1 port map( A => n20015, ZN => n19997);
   U87 : INV_X1 port map( A => n20015, ZN => n19996);
   U88 : INV_X1 port map( A => n20239, ZN => n20222);
   U89 : INV_X1 port map( A => n20239, ZN => n20221);
   U90 : INV_X1 port map( A => n20239, ZN => n20220);
   U91 : INV_X1 port map( A => n19511, ZN => n19492);
   U92 : INV_X1 port map( A => n19511, ZN => n19493);
   U93 : INV_X1 port map( A => n19511, ZN => n19494);
   U94 : INV_X1 port map( A => n19595, ZN => n19578);
   U95 : INV_X1 port map( A => n19595, ZN => n19577);
   U96 : INV_X1 port map( A => n19595, ZN => n19576);
   U97 : INV_X1 port map( A => n19819, ZN => n19802);
   U98 : INV_X1 port map( A => n19819, ZN => n19801);
   U99 : INV_X1 port map( A => n19819, ZN => n19800);
   U100 : INV_X1 port map( A => n19707, ZN => n19690);
   U101 : INV_X1 port map( A => n19707, ZN => n19689);
   U102 : INV_X1 port map( A => n19707, ZN => n19688);
   U103 : INV_X1 port map( A => n19931, ZN => n19914);
   U104 : INV_X1 port map( A => n19931, ZN => n19913);
   U105 : INV_X1 port map( A => n19931, ZN => n19912);
   U106 : INV_X1 port map( A => n20155, ZN => n20138);
   U107 : INV_X1 port map( A => n20155, ZN => n20137);
   U108 : INV_X1 port map( A => n20155, ZN => n20136);
   U109 : INV_X1 port map( A => n20099, ZN => n20082);
   U110 : INV_X1 port map( A => n20099, ZN => n20081);
   U111 : INV_X1 port map( A => n20099, ZN => n20080);
   U112 : INV_X1 port map( A => n19651, ZN => n19634);
   U113 : INV_X1 port map( A => n19651, ZN => n19633);
   U114 : INV_X1 port map( A => n19651, ZN => n19632);
   U115 : INV_X1 port map( A => n20323, ZN => n20306);
   U116 : INV_X1 port map( A => n20323, ZN => n20305);
   U117 : INV_X1 port map( A => n20323, ZN => n20304);
   U118 : INV_X1 port map( A => n19987, ZN => n19970);
   U119 : INV_X1 port map( A => n19987, ZN => n19969);
   U120 : INV_X1 port map( A => n19987, ZN => n19968);
   U121 : INV_X1 port map( A => n20211, ZN => n20194);
   U122 : INV_X1 port map( A => n20211, ZN => n20193);
   U123 : INV_X1 port map( A => n20211, ZN => n20192);
   U124 : INV_X1 port map( A => n19539, ZN => n19522);
   U125 : INV_X1 port map( A => n19539, ZN => n19521);
   U126 : INV_X1 port map( A => n19539, ZN => n19520);
   U127 : INV_X1 port map( A => n19875, ZN => n19858);
   U128 : INV_X1 port map( A => n19875, ZN => n19857);
   U129 : INV_X1 port map( A => n19875, ZN => n19856);
   U130 : INV_X1 port map( A => n19763, ZN => n19746);
   U131 : INV_X1 port map( A => n19763, ZN => n19745);
   U132 : INV_X1 port map( A => n19763, ZN => n19744);
   U133 : INV_X1 port map( A => n20043, ZN => n20026);
   U134 : INV_X1 port map( A => n20043, ZN => n20025);
   U135 : INV_X1 port map( A => n20043, ZN => n20024);
   U136 : INV_X1 port map( A => n20571, ZN => n20554);
   U137 : INV_X1 port map( A => n20571, ZN => n20553);
   U138 : INV_X1 port map( A => n20571, ZN => n20552);
   U139 : INV_X1 port map( A => n20267, ZN => n20250);
   U140 : INV_X1 port map( A => n20267, ZN => n20249);
   U141 : INV_X1 port map( A => n20267, ZN => n20248);
   U142 : BUF_X1 port map( A => n19824, Z => n19845);
   U143 : BUF_X1 port map( A => n19824, Z => n19844);
   U144 : BUF_X1 port map( A => n19824, Z => n19843);
   U145 : BUF_X1 port map( A => n19823, Z => n19842);
   U146 : BUF_X1 port map( A => n19823, Z => n19841);
   U147 : BUF_X1 port map( A => n19823, Z => n19840);
   U148 : BUF_X1 port map( A => n19822, Z => n19839);
   U149 : BUF_X1 port map( A => n19822, Z => n19838);
   U150 : BUF_X1 port map( A => n19822, Z => n19837);
   U151 : BUF_X1 port map( A => n19821, Z => n19836);
   U152 : BUF_X1 port map( A => n19821, Z => n19835);
   U153 : BUF_X1 port map( A => n19821, Z => n19834);
   U154 : BUF_X1 port map( A => n19820, Z => n19833);
   U155 : BUF_X1 port map( A => n19820, Z => n19832);
   U156 : BUF_X1 port map( A => n19820, Z => n19831);
   U157 : BUF_X1 port map( A => n19712, Z => n19733);
   U158 : BUF_X1 port map( A => n19712, Z => n19732);
   U159 : BUF_X1 port map( A => n19712, Z => n19731);
   U160 : BUF_X1 port map( A => n19711, Z => n19730);
   U161 : BUF_X1 port map( A => n19711, Z => n19729);
   U162 : BUF_X1 port map( A => n19711, Z => n19728);
   U163 : BUF_X1 port map( A => n19710, Z => n19727);
   U164 : BUF_X1 port map( A => n19710, Z => n19726);
   U165 : BUF_X1 port map( A => n19710, Z => n19725);
   U166 : BUF_X1 port map( A => n19709, Z => n19724);
   U167 : BUF_X1 port map( A => n19709, Z => n19723);
   U168 : BUF_X1 port map( A => n19709, Z => n19722);
   U169 : BUF_X1 port map( A => n19708, Z => n19721);
   U170 : BUF_X1 port map( A => n19708, Z => n19720);
   U171 : BUF_X1 port map( A => n19708, Z => n19719);
   U172 : BUF_X1 port map( A => n20048, Z => n20069);
   U173 : BUF_X1 port map( A => n20048, Z => n20068);
   U174 : BUF_X1 port map( A => n20048, Z => n20067);
   U175 : BUF_X1 port map( A => n20047, Z => n20066);
   U176 : BUF_X1 port map( A => n20047, Z => n20065);
   U177 : BUF_X1 port map( A => n20047, Z => n20064);
   U178 : BUF_X1 port map( A => n20046, Z => n20063);
   U179 : BUF_X1 port map( A => n20046, Z => n20062);
   U180 : BUF_X1 port map( A => n20046, Z => n20061);
   U181 : BUF_X1 port map( A => n20045, Z => n20060);
   U182 : BUF_X1 port map( A => n20045, Z => n20059);
   U183 : BUF_X1 port map( A => n20045, Z => n20058);
   U184 : BUF_X1 port map( A => n20044, Z => n20057);
   U185 : BUF_X1 port map( A => n20044, Z => n20056);
   U186 : BUF_X1 port map( A => n20044, Z => n20055);
   U187 : BUF_X1 port map( A => n19656, Z => n19677);
   U188 : BUF_X1 port map( A => n19656, Z => n19676);
   U189 : BUF_X1 port map( A => n19656, Z => n19675);
   U190 : BUF_X1 port map( A => n19655, Z => n19674);
   U191 : BUF_X1 port map( A => n19655, Z => n19673);
   U192 : BUF_X1 port map( A => n19655, Z => n19672);
   U193 : BUF_X1 port map( A => n19654, Z => n19671);
   U194 : BUF_X1 port map( A => n19654, Z => n19670);
   U195 : BUF_X1 port map( A => n19654, Z => n19669);
   U196 : BUF_X1 port map( A => n19653, Z => n19668);
   U197 : BUF_X1 port map( A => n19653, Z => n19667);
   U198 : BUF_X1 port map( A => n19653, Z => n19666);
   U199 : BUF_X1 port map( A => n19652, Z => n19665);
   U200 : BUF_X1 port map( A => n19652, Z => n19664);
   U201 : BUF_X1 port map( A => n19652, Z => n19663);
   U202 : BUF_X1 port map( A => n20272, Z => n20293);
   U203 : BUF_X1 port map( A => n20272, Z => n20292);
   U204 : BUF_X1 port map( A => n20272, Z => n20291);
   U205 : BUF_X1 port map( A => n20271, Z => n20290);
   U206 : BUF_X1 port map( A => n20271, Z => n20289);
   U207 : BUF_X1 port map( A => n20271, Z => n20288);
   U208 : BUF_X1 port map( A => n20270, Z => n20287);
   U209 : BUF_X1 port map( A => n20270, Z => n20286);
   U210 : BUF_X1 port map( A => n20270, Z => n20285);
   U211 : BUF_X1 port map( A => n20269, Z => n20284);
   U212 : BUF_X1 port map( A => n20269, Z => n20283);
   U213 : BUF_X1 port map( A => n20269, Z => n20282);
   U214 : BUF_X1 port map( A => n20268, Z => n20281);
   U215 : BUF_X1 port map( A => n20268, Z => n20280);
   U216 : BUF_X1 port map( A => n20268, Z => n20279);
   U217 : BUF_X1 port map( A => n19936, Z => n19957);
   U218 : BUF_X1 port map( A => n19936, Z => n19956);
   U219 : BUF_X1 port map( A => n19936, Z => n19955);
   U220 : BUF_X1 port map( A => n19935, Z => n19954);
   U221 : BUF_X1 port map( A => n19935, Z => n19953);
   U222 : BUF_X1 port map( A => n19935, Z => n19952);
   U223 : BUF_X1 port map( A => n19934, Z => n19951);
   U224 : BUF_X1 port map( A => n19934, Z => n19950);
   U225 : BUF_X1 port map( A => n19934, Z => n19949);
   U226 : BUF_X1 port map( A => n19933, Z => n19948);
   U227 : BUF_X1 port map( A => n19933, Z => n19947);
   U228 : BUF_X1 port map( A => n19933, Z => n19946);
   U229 : BUF_X1 port map( A => n19932, Z => n19945);
   U230 : BUF_X1 port map( A => n19932, Z => n19944);
   U231 : BUF_X1 port map( A => n19932, Z => n19943);
   U232 : BUF_X1 port map( A => n20160, Z => n20181);
   U233 : BUF_X1 port map( A => n20160, Z => n20180);
   U234 : BUF_X1 port map( A => n20160, Z => n20179);
   U235 : BUF_X1 port map( A => n20159, Z => n20178);
   U236 : BUF_X1 port map( A => n20159, Z => n20177);
   U237 : BUF_X1 port map( A => n20159, Z => n20176);
   U238 : BUF_X1 port map( A => n20158, Z => n20175);
   U239 : BUF_X1 port map( A => n20158, Z => n20174);
   U240 : BUF_X1 port map( A => n20158, Z => n20173);
   U241 : BUF_X1 port map( A => n20157, Z => n20172);
   U242 : BUF_X1 port map( A => n20157, Z => n20171);
   U243 : BUF_X1 port map( A => n20157, Z => n20170);
   U244 : BUF_X1 port map( A => n20156, Z => n20169);
   U245 : BUF_X1 port map( A => n20156, Z => n20168);
   U246 : BUF_X1 port map( A => n20156, Z => n20167);
   U247 : BUF_X1 port map( A => n19768, Z => n19789);
   U248 : BUF_X1 port map( A => n19768, Z => n19788);
   U249 : BUF_X1 port map( A => n19768, Z => n19787);
   U250 : BUF_X1 port map( A => n19767, Z => n19786);
   U251 : BUF_X1 port map( A => n19767, Z => n19785);
   U252 : BUF_X1 port map( A => n19767, Z => n19784);
   U253 : BUF_X1 port map( A => n19766, Z => n19783);
   U254 : BUF_X1 port map( A => n19766, Z => n19782);
   U255 : BUF_X1 port map( A => n19766, Z => n19781);
   U256 : BUF_X1 port map( A => n19765, Z => n19780);
   U257 : BUF_X1 port map( A => n19765, Z => n19779);
   U258 : BUF_X1 port map( A => n19765, Z => n19778);
   U259 : BUF_X1 port map( A => n19764, Z => n19777);
   U260 : BUF_X1 port map( A => n19764, Z => n19776);
   U261 : BUF_X1 port map( A => n19764, Z => n19775);
   U262 : BUF_X1 port map( A => n20328, Z => n20349);
   U263 : BUF_X1 port map( A => n20328, Z => n20348);
   U264 : BUF_X1 port map( A => n20328, Z => n20347);
   U265 : BUF_X1 port map( A => n20327, Z => n20346);
   U266 : BUF_X1 port map( A => n20327, Z => n20345);
   U267 : BUF_X1 port map( A => n20327, Z => n20344);
   U268 : BUF_X1 port map( A => n20326, Z => n20343);
   U269 : BUF_X1 port map( A => n20326, Z => n20342);
   U270 : BUF_X1 port map( A => n20326, Z => n20341);
   U271 : BUF_X1 port map( A => n20325, Z => n20340);
   U272 : BUF_X1 port map( A => n20325, Z => n20339);
   U273 : BUF_X1 port map( A => n20325, Z => n20338);
   U274 : BUF_X1 port map( A => n20324, Z => n20337);
   U275 : BUF_X1 port map( A => n20324, Z => n20336);
   U276 : BUF_X1 port map( A => n20324, Z => n20335);
   U277 : BUF_X1 port map( A => n20216, Z => n20237);
   U278 : BUF_X1 port map( A => n20216, Z => n20236);
   U279 : BUF_X1 port map( A => n20216, Z => n20235);
   U280 : BUF_X1 port map( A => n20215, Z => n20234);
   U281 : BUF_X1 port map( A => n20215, Z => n20233);
   U282 : BUF_X1 port map( A => n20215, Z => n20232);
   U283 : BUF_X1 port map( A => n20214, Z => n20231);
   U284 : BUF_X1 port map( A => n20214, Z => n20230);
   U285 : BUF_X1 port map( A => n20214, Z => n20229);
   U286 : BUF_X1 port map( A => n20213, Z => n20228);
   U287 : BUF_X1 port map( A => n20213, Z => n20227);
   U288 : BUF_X1 port map( A => n20213, Z => n20226);
   U289 : BUF_X1 port map( A => n20212, Z => n20225);
   U290 : BUF_X1 port map( A => n20212, Z => n20224);
   U291 : BUF_X1 port map( A => n20212, Z => n20223);
   U292 : BUF_X1 port map( A => n19825, Z => n19846);
   U293 : BUF_X1 port map( A => n19713, Z => n19734);
   U294 : BUF_X1 port map( A => n20049, Z => n20070);
   U295 : BUF_X1 port map( A => n19657, Z => n19678);
   U296 : BUF_X1 port map( A => n20273, Z => n20294);
   U297 : BUF_X1 port map( A => n19937, Z => n19958);
   U298 : BUF_X1 port map( A => n20161, Z => n20182);
   U299 : BUF_X1 port map( A => n19769, Z => n19790);
   U300 : BUF_X1 port map( A => n20329, Z => n20350);
   U301 : BUF_X1 port map( A => n20217, Z => n20238);
   U302 : BUF_X1 port map( A => n19600, Z => n19621);
   U303 : BUF_X1 port map( A => n19600, Z => n19620);
   U304 : BUF_X1 port map( A => n19600, Z => n19619);
   U305 : BUF_X1 port map( A => n19599, Z => n19618);
   U306 : BUF_X1 port map( A => n19599, Z => n19617);
   U307 : BUF_X1 port map( A => n19599, Z => n19616);
   U308 : BUF_X1 port map( A => n19598, Z => n19615);
   U309 : BUF_X1 port map( A => n19598, Z => n19614);
   U310 : BUF_X1 port map( A => n19598, Z => n19613);
   U311 : BUF_X1 port map( A => n19597, Z => n19612);
   U312 : BUF_X1 port map( A => n19597, Z => n19611);
   U313 : BUF_X1 port map( A => n19597, Z => n19610);
   U314 : BUF_X1 port map( A => n19596, Z => n19609);
   U315 : BUF_X1 port map( A => n19596, Z => n19608);
   U316 : BUF_X1 port map( A => n19596, Z => n19607);
   U317 : BUF_X1 port map( A => n20104, Z => n20125);
   U318 : BUF_X1 port map( A => n20104, Z => n20124);
   U319 : BUF_X1 port map( A => n20104, Z => n20123);
   U320 : BUF_X1 port map( A => n20103, Z => n20122);
   U321 : BUF_X1 port map( A => n20103, Z => n20121);
   U322 : BUF_X1 port map( A => n20103, Z => n20120);
   U323 : BUF_X1 port map( A => n20102, Z => n20119);
   U324 : BUF_X1 port map( A => n20102, Z => n20118);
   U325 : BUF_X1 port map( A => n20102, Z => n20117);
   U326 : BUF_X1 port map( A => n20101, Z => n20116);
   U327 : BUF_X1 port map( A => n20101, Z => n20115);
   U328 : BUF_X1 port map( A => n20101, Z => n20114);
   U329 : BUF_X1 port map( A => n20100, Z => n20113);
   U330 : BUF_X1 port map( A => n20100, Z => n20112);
   U331 : BUF_X1 port map( A => n20100, Z => n20111);
   U332 : BUF_X1 port map( A => n19880, Z => n19901);
   U333 : BUF_X1 port map( A => n19880, Z => n19900);
   U334 : BUF_X1 port map( A => n19880, Z => n19899);
   U335 : BUF_X1 port map( A => n19879, Z => n19898);
   U336 : BUF_X1 port map( A => n19879, Z => n19897);
   U337 : BUF_X1 port map( A => n19879, Z => n19896);
   U338 : BUF_X1 port map( A => n19878, Z => n19895);
   U339 : BUF_X1 port map( A => n19878, Z => n19894);
   U340 : BUF_X1 port map( A => n19878, Z => n19893);
   U341 : BUF_X1 port map( A => n19877, Z => n19892);
   U342 : BUF_X1 port map( A => n19877, Z => n19891);
   U343 : BUF_X1 port map( A => n19877, Z => n19890);
   U344 : BUF_X1 port map( A => n19876, Z => n19889);
   U345 : BUF_X1 port map( A => n19876, Z => n19888);
   U346 : BUF_X1 port map( A => n19876, Z => n19887);
   U347 : BUF_X1 port map( A => n19544, Z => n19565);
   U348 : BUF_X1 port map( A => n19544, Z => n19564);
   U349 : BUF_X1 port map( A => n19544, Z => n19563);
   U350 : BUF_X1 port map( A => n19543, Z => n19562);
   U351 : BUF_X1 port map( A => n19543, Z => n19561);
   U352 : BUF_X1 port map( A => n19543, Z => n19560);
   U353 : BUF_X1 port map( A => n19542, Z => n19559);
   U354 : BUF_X1 port map( A => n19542, Z => n19558);
   U355 : BUF_X1 port map( A => n19542, Z => n19557);
   U356 : BUF_X1 port map( A => n19541, Z => n19556);
   U357 : BUF_X1 port map( A => n19541, Z => n19555);
   U358 : BUF_X1 port map( A => n19541, Z => n19554);
   U359 : BUF_X1 port map( A => n19540, Z => n19553);
   U360 : BUF_X1 port map( A => n19540, Z => n19552);
   U361 : BUF_X1 port map( A => n19540, Z => n19551);
   U362 : BUF_X1 port map( A => n19992, Z => n20013);
   U363 : BUF_X1 port map( A => n19992, Z => n20012);
   U364 : BUF_X1 port map( A => n19992, Z => n20011);
   U365 : BUF_X1 port map( A => n19991, Z => n20010);
   U366 : BUF_X1 port map( A => n19991, Z => n20009);
   U367 : BUF_X1 port map( A => n19991, Z => n20008);
   U368 : BUF_X1 port map( A => n19990, Z => n20007);
   U369 : BUF_X1 port map( A => n19990, Z => n20006);
   U370 : BUF_X1 port map( A => n19990, Z => n20005);
   U371 : BUF_X1 port map( A => n19989, Z => n20004);
   U372 : BUF_X1 port map( A => n19989, Z => n20003);
   U373 : BUF_X1 port map( A => n19989, Z => n20002);
   U374 : BUF_X1 port map( A => n19988, Z => n20001);
   U375 : BUF_X1 port map( A => n19988, Z => n20000);
   U376 : BUF_X1 port map( A => n19988, Z => n19999);
   U377 : BUF_X1 port map( A => n19601, Z => n19622);
   U378 : BUF_X1 port map( A => n20105, Z => n20126);
   U379 : BUF_X1 port map( A => n19881, Z => n19902);
   U380 : BUF_X1 port map( A => n19545, Z => n19566);
   U381 : BUF_X1 port map( A => n19993, Z => n20014);
   U382 : BUF_X1 port map( A => n19484, Z => n19495);
   U383 : BUF_X1 port map( A => n19488, Z => n19507);
   U384 : BUF_X1 port map( A => n19487, Z => n19506);
   U385 : BUF_X1 port map( A => n19487, Z => n19505);
   U386 : BUF_X1 port map( A => n19487, Z => n19504);
   U387 : BUF_X1 port map( A => n19486, Z => n19502);
   U388 : BUF_X1 port map( A => n19486, Z => n19501);
   U389 : BUF_X1 port map( A => n19485, Z => n19500);
   U390 : BUF_X1 port map( A => n19485, Z => n19499);
   U391 : BUF_X1 port map( A => n19485, Z => n19498);
   U392 : BUF_X1 port map( A => n19484, Z => n19497);
   U393 : BUF_X1 port map( A => n19488, Z => n19509);
   U394 : BUF_X1 port map( A => n19488, Z => n19508);
   U395 : BUF_X1 port map( A => n19484, Z => n19496);
   U396 : BUF_X1 port map( A => n19486, Z => n19503);
   U397 : BUF_X1 port map( A => n19489, Z => n19510);
   U398 : BUF_X1 port map( A => n3158, Z => n19018);
   U399 : BUF_X1 port map( A => n3158, Z => n19015);
   U400 : BUF_X1 port map( A => n3158, Z => n19016);
   U401 : BUF_X1 port map( A => n3158, Z => n19017);
   U402 : BUF_X1 port map( A => n3114, Z => n19183);
   U403 : BUF_X1 port map( A => n2995, Z => n19382);
   U404 : BUF_X1 port map( A => n3114, Z => n19184);
   U405 : BUF_X1 port map( A => n2995, Z => n19383);
   U406 : BUF_X1 port map( A => n3114, Z => n19185);
   U407 : BUF_X1 port map( A => n2995, Z => n19384);
   U408 : BUF_X1 port map( A => n3114, Z => n19186);
   U409 : BUF_X1 port map( A => n2995, Z => n19385);
   U410 : BUF_X1 port map( A => n3114, Z => n19187);
   U411 : BUF_X1 port map( A => n2995, Z => n19386);
   U412 : BUF_X1 port map( A => n3135, Z => n19086);
   U413 : BUF_X1 port map( A => n3135, Z => n19087);
   U414 : BUF_X1 port map( A => n3135, Z => n19088);
   U415 : BUF_X1 port map( A => n3135, Z => n19089);
   U416 : BUF_X1 port map( A => n3135, Z => n19090);
   U417 : BUF_X1 port map( A => n3019, Z => n19285);
   U418 : BUF_X1 port map( A => n3019, Z => n19286);
   U419 : BUF_X1 port map( A => n3019, Z => n19287);
   U420 : BUF_X1 port map( A => n3019, Z => n19288);
   U421 : BUF_X1 port map( A => n3019, Z => n19289);
   U422 : BUF_X1 port map( A => n19165, Z => n19170);
   U423 : BUF_X1 port map( A => n19364, Z => n19369);
   U424 : BUF_X1 port map( A => n19165, Z => n19169);
   U425 : BUF_X1 port map( A => n19364, Z => n19368);
   U426 : BUF_X1 port map( A => n19164, Z => n19168);
   U427 : BUF_X1 port map( A => n19363, Z => n19367);
   U428 : BUF_X1 port map( A => n19164, Z => n19167);
   U429 : BUF_X1 port map( A => n19363, Z => n19366);
   U430 : BUF_X1 port map( A => n3122, Z => n19158);
   U431 : BUF_X1 port map( A => n3005, Z => n19357);
   U432 : BUF_X1 port map( A => n3122, Z => n19159);
   U433 : BUF_X1 port map( A => n3005, Z => n19358);
   U434 : BUF_X1 port map( A => n3122, Z => n19160);
   U435 : BUF_X1 port map( A => n3005, Z => n19359);
   U436 : BUF_X1 port map( A => n3122, Z => n19161);
   U437 : BUF_X1 port map( A => n3005, Z => n19360);
   U438 : BUF_X1 port map( A => n3122, Z => n19162);
   U439 : BUF_X1 port map( A => n3005, Z => n19361);
   U440 : BUF_X1 port map( A => n3112, Z => n19189);
   U441 : BUF_X1 port map( A => n2993, Z => n19388);
   U442 : BUF_X1 port map( A => n3112, Z => n19190);
   U443 : BUF_X1 port map( A => n2993, Z => n19389);
   U444 : BUF_X1 port map( A => n3112, Z => n19191);
   U445 : BUF_X1 port map( A => n2993, Z => n19390);
   U446 : BUF_X1 port map( A => n3112, Z => n19192);
   U447 : BUF_X1 port map( A => n2993, Z => n19391);
   U448 : BUF_X1 port map( A => n3112, Z => n19193);
   U449 : BUF_X1 port map( A => n2993, Z => n19392);
   U450 : BUF_X1 port map( A => n19164, Z => n19166);
   U451 : BUF_X1 port map( A => n19363, Z => n19365);
   U452 : BUF_X1 port map( A => n3158, Z => n19014);
   U453 : BUF_X1 port map( A => n19684, Z => n19705);
   U454 : BUF_X1 port map( A => n19684, Z => n19704);
   U455 : BUF_X1 port map( A => n19684, Z => n19703);
   U456 : BUF_X1 port map( A => n19683, Z => n19702);
   U457 : BUF_X1 port map( A => n19683, Z => n19701);
   U458 : BUF_X1 port map( A => n19683, Z => n19700);
   U459 : BUF_X1 port map( A => n19682, Z => n19699);
   U460 : BUF_X1 port map( A => n19682, Z => n19698);
   U461 : BUF_X1 port map( A => n19682, Z => n19697);
   U462 : BUF_X1 port map( A => n19681, Z => n19696);
   U463 : BUF_X1 port map( A => n19681, Z => n19695);
   U464 : BUF_X1 port map( A => n19681, Z => n19694);
   U465 : BUF_X1 port map( A => n19680, Z => n19693);
   U466 : BUF_X1 port map( A => n19680, Z => n19692);
   U467 : BUF_X1 port map( A => n19680, Z => n19691);
   U468 : BUF_X1 port map( A => n20132, Z => n20153);
   U469 : BUF_X1 port map( A => n20132, Z => n20152);
   U470 : BUF_X1 port map( A => n20132, Z => n20151);
   U471 : BUF_X1 port map( A => n20131, Z => n20150);
   U472 : BUF_X1 port map( A => n20131, Z => n20149);
   U473 : BUF_X1 port map( A => n20131, Z => n20148);
   U474 : BUF_X1 port map( A => n20130, Z => n20147);
   U475 : BUF_X1 port map( A => n20130, Z => n20146);
   U476 : BUF_X1 port map( A => n20130, Z => n20145);
   U477 : BUF_X1 port map( A => n20129, Z => n20144);
   U478 : BUF_X1 port map( A => n20129, Z => n20143);
   U479 : BUF_X1 port map( A => n20129, Z => n20142);
   U480 : BUF_X1 port map( A => n20128, Z => n20141);
   U481 : BUF_X1 port map( A => n20128, Z => n20140);
   U482 : BUF_X1 port map( A => n20128, Z => n20139);
   U483 : BUF_X1 port map( A => n19628, Z => n19649);
   U484 : BUF_X1 port map( A => n19628, Z => n19648);
   U485 : BUF_X1 port map( A => n19628, Z => n19647);
   U486 : BUF_X1 port map( A => n19627, Z => n19646);
   U487 : BUF_X1 port map( A => n19627, Z => n19645);
   U488 : BUF_X1 port map( A => n19627, Z => n19644);
   U489 : BUF_X1 port map( A => n19626, Z => n19643);
   U490 : BUF_X1 port map( A => n19626, Z => n19642);
   U491 : BUF_X1 port map( A => n19626, Z => n19641);
   U492 : BUF_X1 port map( A => n19625, Z => n19640);
   U493 : BUF_X1 port map( A => n19625, Z => n19639);
   U494 : BUF_X1 port map( A => n19625, Z => n19638);
   U495 : BUF_X1 port map( A => n19624, Z => n19637);
   U496 : BUF_X1 port map( A => n19624, Z => n19636);
   U497 : BUF_X1 port map( A => n19624, Z => n19635);
   U498 : BUF_X1 port map( A => n20300, Z => n20321);
   U499 : BUF_X1 port map( A => n20300, Z => n20320);
   U500 : BUF_X1 port map( A => n20300, Z => n20319);
   U501 : BUF_X1 port map( A => n20299, Z => n20318);
   U502 : BUF_X1 port map( A => n20299, Z => n20317);
   U503 : BUF_X1 port map( A => n20299, Z => n20316);
   U504 : BUF_X1 port map( A => n20298, Z => n20315);
   U505 : BUF_X1 port map( A => n20298, Z => n20314);
   U506 : BUF_X1 port map( A => n20298, Z => n20313);
   U507 : BUF_X1 port map( A => n20297, Z => n20312);
   U508 : BUF_X1 port map( A => n20297, Z => n20311);
   U509 : BUF_X1 port map( A => n20297, Z => n20310);
   U510 : BUF_X1 port map( A => n20296, Z => n20309);
   U511 : BUF_X1 port map( A => n20296, Z => n20308);
   U512 : BUF_X1 port map( A => n20296, Z => n20307);
   U513 : BUF_X1 port map( A => n19964, Z => n19985);
   U514 : BUF_X1 port map( A => n19964, Z => n19984);
   U515 : BUF_X1 port map( A => n19964, Z => n19983);
   U516 : BUF_X1 port map( A => n19963, Z => n19982);
   U517 : BUF_X1 port map( A => n19963, Z => n19981);
   U518 : BUF_X1 port map( A => n19963, Z => n19980);
   U519 : BUF_X1 port map( A => n19962, Z => n19979);
   U520 : BUF_X1 port map( A => n19962, Z => n19978);
   U521 : BUF_X1 port map( A => n19962, Z => n19977);
   U522 : BUF_X1 port map( A => n19961, Z => n19976);
   U523 : BUF_X1 port map( A => n19961, Z => n19975);
   U524 : BUF_X1 port map( A => n19961, Z => n19974);
   U525 : BUF_X1 port map( A => n19960, Z => n19973);
   U526 : BUF_X1 port map( A => n19960, Z => n19972);
   U527 : BUF_X1 port map( A => n19960, Z => n19971);
   U528 : BUF_X1 port map( A => n20188, Z => n20209);
   U529 : BUF_X1 port map( A => n20188, Z => n20208);
   U530 : BUF_X1 port map( A => n20188, Z => n20207);
   U531 : BUF_X1 port map( A => n20187, Z => n20206);
   U532 : BUF_X1 port map( A => n20187, Z => n20205);
   U533 : BUF_X1 port map( A => n20187, Z => n20204);
   U534 : BUF_X1 port map( A => n20186, Z => n20203);
   U535 : BUF_X1 port map( A => n20186, Z => n20202);
   U536 : BUF_X1 port map( A => n20186, Z => n20201);
   U537 : BUF_X1 port map( A => n20185, Z => n20200);
   U538 : BUF_X1 port map( A => n20185, Z => n20199);
   U539 : BUF_X1 port map( A => n20185, Z => n20198);
   U540 : BUF_X1 port map( A => n20184, Z => n20197);
   U541 : BUF_X1 port map( A => n20184, Z => n20196);
   U542 : BUF_X1 port map( A => n20184, Z => n20195);
   U543 : BUF_X1 port map( A => n19516, Z => n19537);
   U544 : BUF_X1 port map( A => n19516, Z => n19536);
   U545 : BUF_X1 port map( A => n19516, Z => n19535);
   U546 : BUF_X1 port map( A => n19515, Z => n19534);
   U547 : BUF_X1 port map( A => n19515, Z => n19533);
   U548 : BUF_X1 port map( A => n19515, Z => n19532);
   U549 : BUF_X1 port map( A => n19514, Z => n19531);
   U550 : BUF_X1 port map( A => n19514, Z => n19530);
   U551 : BUF_X1 port map( A => n19514, Z => n19529);
   U552 : BUF_X1 port map( A => n19513, Z => n19528);
   U553 : BUF_X1 port map( A => n19513, Z => n19527);
   U554 : BUF_X1 port map( A => n19513, Z => n19526);
   U555 : BUF_X1 port map( A => n19512, Z => n19525);
   U556 : BUF_X1 port map( A => n19512, Z => n19524);
   U557 : BUF_X1 port map( A => n19512, Z => n19523);
   U558 : BUF_X1 port map( A => n19852, Z => n19873);
   U559 : BUF_X1 port map( A => n19852, Z => n19872);
   U560 : BUF_X1 port map( A => n19852, Z => n19871);
   U561 : BUF_X1 port map( A => n19851, Z => n19870);
   U562 : BUF_X1 port map( A => n19851, Z => n19869);
   U563 : BUF_X1 port map( A => n19851, Z => n19868);
   U564 : BUF_X1 port map( A => n19850, Z => n19867);
   U565 : BUF_X1 port map( A => n19850, Z => n19866);
   U566 : BUF_X1 port map( A => n19850, Z => n19865);
   U567 : BUF_X1 port map( A => n19849, Z => n19864);
   U568 : BUF_X1 port map( A => n19849, Z => n19863);
   U569 : BUF_X1 port map( A => n19849, Z => n19862);
   U570 : BUF_X1 port map( A => n19848, Z => n19861);
   U571 : BUF_X1 port map( A => n19848, Z => n19860);
   U572 : BUF_X1 port map( A => n19848, Z => n19859);
   U573 : BUF_X1 port map( A => n19740, Z => n19761);
   U574 : BUF_X1 port map( A => n19740, Z => n19760);
   U575 : BUF_X1 port map( A => n19740, Z => n19759);
   U576 : BUF_X1 port map( A => n19739, Z => n19758);
   U577 : BUF_X1 port map( A => n19739, Z => n19757);
   U578 : BUF_X1 port map( A => n19739, Z => n19756);
   U579 : BUF_X1 port map( A => n19738, Z => n19755);
   U580 : BUF_X1 port map( A => n19738, Z => n19754);
   U581 : BUF_X1 port map( A => n19738, Z => n19753);
   U582 : BUF_X1 port map( A => n19737, Z => n19752);
   U583 : BUF_X1 port map( A => n19737, Z => n19751);
   U584 : BUF_X1 port map( A => n19737, Z => n19750);
   U585 : BUF_X1 port map( A => n19736, Z => n19749);
   U586 : BUF_X1 port map( A => n19736, Z => n19748);
   U587 : BUF_X1 port map( A => n19736, Z => n19747);
   U588 : BUF_X1 port map( A => n20020, Z => n20041);
   U589 : BUF_X1 port map( A => n20020, Z => n20040);
   U590 : BUF_X1 port map( A => n20020, Z => n20039);
   U591 : BUF_X1 port map( A => n20019, Z => n20038);
   U592 : BUF_X1 port map( A => n20019, Z => n20037);
   U593 : BUF_X1 port map( A => n20019, Z => n20036);
   U594 : BUF_X1 port map( A => n20018, Z => n20035);
   U595 : BUF_X1 port map( A => n20018, Z => n20034);
   U596 : BUF_X1 port map( A => n20018, Z => n20033);
   U597 : BUF_X1 port map( A => n20017, Z => n20032);
   U598 : BUF_X1 port map( A => n20017, Z => n20031);
   U599 : BUF_X1 port map( A => n20017, Z => n20030);
   U600 : BUF_X1 port map( A => n20016, Z => n20029);
   U601 : BUF_X1 port map( A => n20016, Z => n20028);
   U602 : BUF_X1 port map( A => n20016, Z => n20027);
   U603 : BUF_X1 port map( A => n20548, Z => n20569);
   U604 : BUF_X1 port map( A => n20548, Z => n20568);
   U605 : BUF_X1 port map( A => n20548, Z => n20567);
   U606 : BUF_X1 port map( A => n20547, Z => n20566);
   U607 : BUF_X1 port map( A => n20547, Z => n20565);
   U608 : BUF_X1 port map( A => n20547, Z => n20564);
   U609 : BUF_X1 port map( A => n20546, Z => n20563);
   U610 : BUF_X1 port map( A => n20546, Z => n20562);
   U611 : BUF_X1 port map( A => n20546, Z => n20561);
   U612 : BUF_X1 port map( A => n20545, Z => n20560);
   U613 : BUF_X1 port map( A => n20545, Z => n20559);
   U614 : BUF_X1 port map( A => n20545, Z => n20558);
   U615 : BUF_X1 port map( A => n20544, Z => n20557);
   U616 : BUF_X1 port map( A => n20544, Z => n20556);
   U617 : BUF_X1 port map( A => n20544, Z => n20555);
   U618 : BUF_X1 port map( A => n20244, Z => n20265);
   U619 : BUF_X1 port map( A => n20244, Z => n20264);
   U620 : BUF_X1 port map( A => n20244, Z => n20263);
   U621 : BUF_X1 port map( A => n20243, Z => n20262);
   U622 : BUF_X1 port map( A => n20243, Z => n20261);
   U623 : BUF_X1 port map( A => n20243, Z => n20260);
   U624 : BUF_X1 port map( A => n20242, Z => n20259);
   U625 : BUF_X1 port map( A => n20242, Z => n20258);
   U626 : BUF_X1 port map( A => n20242, Z => n20257);
   U627 : BUF_X1 port map( A => n20241, Z => n20256);
   U628 : BUF_X1 port map( A => n20241, Z => n20255);
   U629 : BUF_X1 port map( A => n20241, Z => n20254);
   U630 : BUF_X1 port map( A => n20240, Z => n20253);
   U631 : BUF_X1 port map( A => n20240, Z => n20252);
   U632 : BUF_X1 port map( A => n20240, Z => n20251);
   U633 : BUF_X1 port map( A => n19685, Z => n19706);
   U634 : BUF_X1 port map( A => n20133, Z => n20154);
   U635 : BUF_X1 port map( A => n19629, Z => n19650);
   U636 : BUF_X1 port map( A => n20301, Z => n20322);
   U637 : BUF_X1 port map( A => n19965, Z => n19986);
   U638 : BUF_X1 port map( A => n20189, Z => n20210);
   U639 : BUF_X1 port map( A => n19517, Z => n19538);
   U640 : BUF_X1 port map( A => n19741, Z => n19762);
   U641 : BUF_X1 port map( A => n19853, Z => n19874);
   U642 : BUF_X1 port map( A => n20021, Z => n20042);
   U643 : BUF_X1 port map( A => n20549, Z => n20570);
   U644 : BUF_X1 port map( A => n20245, Z => n20266);
   U645 : BUF_X1 port map( A => n19572, Z => n19593);
   U646 : BUF_X1 port map( A => n19572, Z => n19592);
   U647 : BUF_X1 port map( A => n19572, Z => n19591);
   U648 : BUF_X1 port map( A => n19571, Z => n19590);
   U649 : BUF_X1 port map( A => n19571, Z => n19589);
   U650 : BUF_X1 port map( A => n19571, Z => n19588);
   U651 : BUF_X1 port map( A => n19570, Z => n19587);
   U652 : BUF_X1 port map( A => n19570, Z => n19586);
   U653 : BUF_X1 port map( A => n19570, Z => n19585);
   U654 : BUF_X1 port map( A => n19569, Z => n19584);
   U655 : BUF_X1 port map( A => n19569, Z => n19583);
   U656 : BUF_X1 port map( A => n19569, Z => n19582);
   U657 : BUF_X1 port map( A => n19568, Z => n19581);
   U658 : BUF_X1 port map( A => n19568, Z => n19580);
   U659 : BUF_X1 port map( A => n19568, Z => n19579);
   U660 : BUF_X1 port map( A => n19796, Z => n19817);
   U661 : BUF_X1 port map( A => n19796, Z => n19816);
   U662 : BUF_X1 port map( A => n19796, Z => n19815);
   U663 : BUF_X1 port map( A => n19795, Z => n19814);
   U664 : BUF_X1 port map( A => n19795, Z => n19813);
   U665 : BUF_X1 port map( A => n19795, Z => n19812);
   U666 : BUF_X1 port map( A => n19794, Z => n19811);
   U667 : BUF_X1 port map( A => n19794, Z => n19810);
   U668 : BUF_X1 port map( A => n19794, Z => n19809);
   U669 : BUF_X1 port map( A => n19793, Z => n19808);
   U670 : BUF_X1 port map( A => n19793, Z => n19807);
   U671 : BUF_X1 port map( A => n19793, Z => n19806);
   U672 : BUF_X1 port map( A => n19792, Z => n19805);
   U673 : BUF_X1 port map( A => n19792, Z => n19804);
   U674 : BUF_X1 port map( A => n19792, Z => n19803);
   U675 : BUF_X1 port map( A => n19908, Z => n19929);
   U676 : BUF_X1 port map( A => n19908, Z => n19928);
   U677 : BUF_X1 port map( A => n19908, Z => n19927);
   U678 : BUF_X1 port map( A => n19907, Z => n19926);
   U679 : BUF_X1 port map( A => n19907, Z => n19925);
   U680 : BUF_X1 port map( A => n19907, Z => n19924);
   U681 : BUF_X1 port map( A => n19906, Z => n19923);
   U682 : BUF_X1 port map( A => n19906, Z => n19922);
   U683 : BUF_X1 port map( A => n19906, Z => n19921);
   U684 : BUF_X1 port map( A => n19905, Z => n19920);
   U685 : BUF_X1 port map( A => n19905, Z => n19919);
   U686 : BUF_X1 port map( A => n19905, Z => n19918);
   U687 : BUF_X1 port map( A => n19904, Z => n19917);
   U688 : BUF_X1 port map( A => n19904, Z => n19916);
   U689 : BUF_X1 port map( A => n19904, Z => n19915);
   U690 : BUF_X1 port map( A => n20076, Z => n20097);
   U691 : BUF_X1 port map( A => n20076, Z => n20096);
   U692 : BUF_X1 port map( A => n20076, Z => n20095);
   U693 : BUF_X1 port map( A => n20075, Z => n20094);
   U694 : BUF_X1 port map( A => n20075, Z => n20093);
   U695 : BUF_X1 port map( A => n20075, Z => n20092);
   U696 : BUF_X1 port map( A => n20074, Z => n20091);
   U697 : BUF_X1 port map( A => n20074, Z => n20090);
   U698 : BUF_X1 port map( A => n20074, Z => n20089);
   U699 : BUF_X1 port map( A => n20073, Z => n20088);
   U700 : BUF_X1 port map( A => n20073, Z => n20087);
   U701 : BUF_X1 port map( A => n20073, Z => n20086);
   U702 : BUF_X1 port map( A => n20072, Z => n20085);
   U703 : BUF_X1 port map( A => n20072, Z => n20084);
   U704 : BUF_X1 port map( A => n20072, Z => n20083);
   U705 : BUF_X1 port map( A => n19573, Z => n19594);
   U706 : BUF_X1 port map( A => n19797, Z => n19818);
   U707 : BUF_X1 port map( A => n19909, Z => n19930);
   U708 : BUF_X1 port map( A => n20077, Z => n20098);
   U709 : BUF_X1 port map( A => n19938, Z => n19936);
   U710 : BUF_X1 port map( A => n19938, Z => n19935);
   U711 : BUF_X1 port map( A => n19939, Z => n19934);
   U712 : BUF_X1 port map( A => n19939, Z => n19933);
   U713 : BUF_X1 port map( A => n19939, Z => n19932);
   U714 : BUF_X1 port map( A => n19658, Z => n19656);
   U715 : BUF_X1 port map( A => n19658, Z => n19655);
   U716 : BUF_X1 port map( A => n19659, Z => n19654);
   U717 : BUF_X1 port map( A => n19659, Z => n19653);
   U718 : BUF_X1 port map( A => n19659, Z => n19652);
   U719 : BUF_X1 port map( A => n19882, Z => n19880);
   U720 : BUF_X1 port map( A => n19882, Z => n19879);
   U721 : BUF_X1 port map( A => n19883, Z => n19878);
   U722 : BUF_X1 port map( A => n19883, Z => n19877);
   U723 : BUF_X1 port map( A => n19883, Z => n19876);
   U724 : BUF_X1 port map( A => n19994, Z => n19992);
   U725 : BUF_X1 port map( A => n19994, Z => n19991);
   U726 : BUF_X1 port map( A => n19995, Z => n19990);
   U727 : BUF_X1 port map( A => n19995, Z => n19989);
   U728 : BUF_X1 port map( A => n19995, Z => n19988);
   U729 : BUF_X1 port map( A => n19770, Z => n19768);
   U730 : BUF_X1 port map( A => n19770, Z => n19767);
   U731 : BUF_X1 port map( A => n19771, Z => n19766);
   U732 : BUF_X1 port map( A => n19771, Z => n19765);
   U733 : BUF_X1 port map( A => n19771, Z => n19764);
   U734 : BUF_X1 port map( A => n19546, Z => n19544);
   U735 : BUF_X1 port map( A => n19546, Z => n19543);
   U736 : BUF_X1 port map( A => n19547, Z => n19542);
   U737 : BUF_X1 port map( A => n19547, Z => n19541);
   U738 : BUF_X1 port map( A => n19547, Z => n19540);
   U739 : BUF_X1 port map( A => n20050, Z => n20048);
   U740 : BUF_X1 port map( A => n20050, Z => n20047);
   U741 : BUF_X1 port map( A => n20051, Z => n20046);
   U742 : BUF_X1 port map( A => n20051, Z => n20045);
   U743 : BUF_X1 port map( A => n20051, Z => n20044);
   U744 : BUF_X1 port map( A => n20106, Z => n20104);
   U745 : BUF_X1 port map( A => n20106, Z => n20103);
   U746 : BUF_X1 port map( A => n20107, Z => n20102);
   U747 : BUF_X1 port map( A => n20107, Z => n20101);
   U748 : BUF_X1 port map( A => n20107, Z => n20100);
   U749 : BUF_X1 port map( A => n20330, Z => n20328);
   U750 : BUF_X1 port map( A => n20330, Z => n20327);
   U751 : BUF_X1 port map( A => n20331, Z => n20326);
   U752 : BUF_X1 port map( A => n20331, Z => n20325);
   U753 : BUF_X1 port map( A => n20331, Z => n20324);
   U754 : BUF_X1 port map( A => n20218, Z => n20216);
   U755 : BUF_X1 port map( A => n20218, Z => n20215);
   U756 : BUF_X1 port map( A => n20219, Z => n20214);
   U757 : BUF_X1 port map( A => n20219, Z => n20213);
   U758 : BUF_X1 port map( A => n20219, Z => n20212);
   U759 : BUF_X1 port map( A => n19826, Z => n19824);
   U760 : BUF_X1 port map( A => n19826, Z => n19823);
   U761 : BUF_X1 port map( A => n19827, Z => n19822);
   U762 : BUF_X1 port map( A => n19827, Z => n19821);
   U763 : BUF_X1 port map( A => n19827, Z => n19820);
   U764 : BUF_X1 port map( A => n19714, Z => n19712);
   U765 : BUF_X1 port map( A => n19714, Z => n19711);
   U766 : BUF_X1 port map( A => n19715, Z => n19710);
   U767 : BUF_X1 port map( A => n19715, Z => n19709);
   U768 : BUF_X1 port map( A => n19715, Z => n19708);
   U769 : BUF_X1 port map( A => n19602, Z => n19600);
   U770 : BUF_X1 port map( A => n19602, Z => n19599);
   U771 : BUF_X1 port map( A => n19603, Z => n19598);
   U772 : BUF_X1 port map( A => n19603, Z => n19597);
   U773 : BUF_X1 port map( A => n19603, Z => n19596);
   U774 : BUF_X1 port map( A => n20274, Z => n20272);
   U775 : BUF_X1 port map( A => n20274, Z => n20271);
   U776 : BUF_X1 port map( A => n20275, Z => n20270);
   U777 : BUF_X1 port map( A => n20275, Z => n20269);
   U778 : BUF_X1 port map( A => n20275, Z => n20268);
   U779 : BUF_X1 port map( A => n20162, Z => n20160);
   U780 : BUF_X1 port map( A => n20162, Z => n20159);
   U781 : BUF_X1 port map( A => n20163, Z => n20158);
   U782 : BUF_X1 port map( A => n20163, Z => n20157);
   U783 : BUF_X1 port map( A => n20163, Z => n20156);
   U784 : BUF_X1 port map( A => n19490, Z => n19487);
   U785 : BUF_X1 port map( A => n19491, Z => n19485);
   U786 : BUF_X1 port map( A => n19490, Z => n19488);
   U787 : BUF_X1 port map( A => n19491, Z => n19484);
   U788 : BUF_X1 port map( A => n19491, Z => n19486);
   U789 : BUF_X1 port map( A => n19938, Z => n19937);
   U790 : BUF_X1 port map( A => n19994, Z => n19993);
   U791 : BUF_X1 port map( A => n19658, Z => n19657);
   U792 : BUF_X1 port map( A => n19882, Z => n19881);
   U793 : BUF_X1 port map( A => n19770, Z => n19769);
   U794 : BUF_X1 port map( A => n19546, Z => n19545);
   U795 : BUF_X1 port map( A => n20050, Z => n20049);
   U796 : BUF_X1 port map( A => n20106, Z => n20105);
   U797 : BUF_X1 port map( A => n20330, Z => n20329);
   U798 : BUF_X1 port map( A => n20218, Z => n20217);
   U799 : BUF_X1 port map( A => n19826, Z => n19825);
   U800 : BUF_X1 port map( A => n19714, Z => n19713);
   U801 : BUF_X1 port map( A => n19602, Z => n19601);
   U802 : BUF_X1 port map( A => n20274, Z => n20273);
   U803 : BUF_X1 port map( A => n20162, Z => n20161);
   U804 : BUF_X1 port map( A => n19490, Z => n19489);
   U805 : NOR2_X1 port map( A1 => n11686, A2 => n11687, ZN => n3158);
   U806 : BUF_X1 port map( A => n3129, Z => n19116);
   U807 : BUF_X1 port map( A => n3129, Z => n19117);
   U808 : BUF_X1 port map( A => n3129, Z => n19118);
   U809 : BUF_X1 port map( A => n3129, Z => n19119);
   U810 : BUF_X1 port map( A => n3129, Z => n19120);
   U811 : BUF_X1 port map( A => n3186, Z => n18940);
   U812 : BUF_X1 port map( A => n3186, Z => n18936);
   U813 : BUF_X1 port map( A => n3186, Z => n18937);
   U814 : BUF_X1 port map( A => n3186, Z => n18938);
   U815 : BUF_X1 port map( A => n3186, Z => n18939);
   U816 : BUF_X1 port map( A => n3134, Z => n19092);
   U817 : BUF_X1 port map( A => n3012, Z => n19315);
   U818 : BUF_X1 port map( A => n3017, Z => n19291);
   U819 : BUF_X1 port map( A => n3134, Z => n19093);
   U820 : BUF_X1 port map( A => n3012, Z => n19316);
   U821 : BUF_X1 port map( A => n3017, Z => n19292);
   U822 : BUF_X1 port map( A => n3134, Z => n19094);
   U823 : BUF_X1 port map( A => n3012, Z => n19317);
   U824 : BUF_X1 port map( A => n3017, Z => n19293);
   U825 : BUF_X1 port map( A => n3134, Z => n19095);
   U826 : BUF_X1 port map( A => n3012, Z => n19318);
   U827 : BUF_X1 port map( A => n3017, Z => n19294);
   U828 : BUF_X1 port map( A => n3134, Z => n19096);
   U829 : BUF_X1 port map( A => n3012, Z => n19319);
   U830 : BUF_X1 port map( A => n3017, Z => n19295);
   U831 : BUF_X1 port map( A => n3109, Z => n19207);
   U832 : BUF_X1 port map( A => n3109, Z => n19208);
   U833 : BUF_X1 port map( A => n3109, Z => n19209);
   U834 : BUF_X1 port map( A => n3109, Z => n19210);
   U835 : BUF_X1 port map( A => n3109, Z => n19211);
   U836 : BUF_X1 port map( A => n3104, Z => n19231);
   U837 : BUF_X1 port map( A => n3035, Z => n19255);
   U838 : BUF_X1 port map( A => n2982, Z => n19430);
   U839 : BUF_X1 port map( A => n2988, Z => n19406);
   U840 : BUF_X1 port map( A => n2783, Z => n19454);
   U841 : BUF_X1 port map( A => n3104, Z => n19232);
   U842 : BUF_X1 port map( A => n3035, Z => n19256);
   U843 : BUF_X1 port map( A => n2982, Z => n19431);
   U844 : BUF_X1 port map( A => n2988, Z => n19407);
   U845 : BUF_X1 port map( A => n2783, Z => n19455);
   U846 : BUF_X1 port map( A => n3104, Z => n19233);
   U847 : BUF_X1 port map( A => n3035, Z => n19257);
   U848 : BUF_X1 port map( A => n2982, Z => n19432);
   U849 : BUF_X1 port map( A => n2988, Z => n19408);
   U850 : BUF_X1 port map( A => n2783, Z => n19456);
   U851 : BUF_X1 port map( A => n3104, Z => n19234);
   U852 : BUF_X1 port map( A => n3035, Z => n19258);
   U853 : BUF_X1 port map( A => n2982, Z => n19433);
   U854 : BUF_X1 port map( A => n2988, Z => n19409);
   U855 : BUF_X1 port map( A => n2783, Z => n19457);
   U856 : BUF_X1 port map( A => n3104, Z => n19235);
   U857 : BUF_X1 port map( A => n3035, Z => n19259);
   U858 : BUF_X1 port map( A => n2982, Z => n19434);
   U859 : BUF_X1 port map( A => n2988, Z => n19410);
   U860 : BUF_X1 port map( A => n2783, Z => n19458);
   U861 : BUF_X1 port map( A => n3130, Z => n19110);
   U862 : BUF_X1 port map( A => n3130, Z => n19111);
   U863 : BUF_X1 port map( A => n3130, Z => n19112);
   U864 : BUF_X1 port map( A => n3130, Z => n19113);
   U865 : BUF_X1 port map( A => n3130, Z => n19114);
   U866 : BUF_X1 port map( A => n3013, Z => n19309);
   U867 : BUF_X1 port map( A => n3013, Z => n19310);
   U868 : BUF_X1 port map( A => n3013, Z => n19311);
   U869 : BUF_X1 port map( A => n3013, Z => n19312);
   U870 : BUF_X1 port map( A => n3013, Z => n19313);
   U871 : BUF_X1 port map( A => n3106, Z => n19220);
   U872 : BUF_X1 port map( A => n3106, Z => n19221);
   U873 : BUF_X1 port map( A => n3106, Z => n19222);
   U874 : BUF_X1 port map( A => n3106, Z => n19223);
   U875 : BUF_X1 port map( A => n2985, Z => n19419);
   U876 : BUF_X1 port map( A => n2985, Z => n19420);
   U877 : BUF_X1 port map( A => n2985, Z => n19421);
   U878 : BUF_X1 port map( A => n2985, Z => n19422);
   U879 : BUF_X1 port map( A => n2780, Z => n19467);
   U880 : BUF_X1 port map( A => n2780, Z => n19468);
   U881 : BUF_X1 port map( A => n2780, Z => n19469);
   U882 : BUF_X1 port map( A => n2780, Z => n19470);
   U883 : BUF_X1 port map( A => n3032, Z => n19268);
   U884 : BUF_X1 port map( A => n3032, Z => n19269);
   U885 : BUF_X1 port map( A => n3032, Z => n19270);
   U886 : BUF_X1 port map( A => n3032, Z => n19271);
   U887 : BUF_X1 port map( A => n3111, Z => n19196);
   U888 : BUF_X1 port map( A => n3037, Z => n19244);
   U889 : BUF_X1 port map( A => n2979, Z => n19443);
   U890 : BUF_X1 port map( A => n2992, Z => n19395);
   U891 : BUF_X1 port map( A => n3111, Z => n19197);
   U892 : BUF_X1 port map( A => n3037, Z => n19245);
   U893 : BUF_X1 port map( A => n2979, Z => n19444);
   U894 : BUF_X1 port map( A => n2992, Z => n19396);
   U895 : BUF_X1 port map( A => n3111, Z => n19198);
   U896 : BUF_X1 port map( A => n3037, Z => n19246);
   U897 : BUF_X1 port map( A => n2979, Z => n19445);
   U898 : BUF_X1 port map( A => n2992, Z => n19397);
   U899 : BUF_X1 port map( A => n3111, Z => n19199);
   U900 : BUF_X1 port map( A => n3037, Z => n19247);
   U901 : BUF_X1 port map( A => n2979, Z => n19446);
   U902 : BUF_X1 port map( A => n2992, Z => n19398);
   U903 : BUF_X1 port map( A => n3128, Z => n19122);
   U904 : BUF_X1 port map( A => n3011, Z => n19321);
   U905 : BUF_X1 port map( A => n3128, Z => n19123);
   U906 : BUF_X1 port map( A => n3011, Z => n19322);
   U907 : BUF_X1 port map( A => n3128, Z => n19124);
   U908 : BUF_X1 port map( A => n3011, Z => n19323);
   U909 : BUF_X1 port map( A => n3128, Z => n19125);
   U910 : BUF_X1 port map( A => n3011, Z => n19324);
   U911 : BUF_X1 port map( A => n3128, Z => n19126);
   U912 : BUF_X1 port map( A => n3011, Z => n19325);
   U913 : BUF_X1 port map( A => n3126, Z => n19134);
   U914 : BUF_X1 port map( A => n3126, Z => n19135);
   U915 : BUF_X1 port map( A => n3126, Z => n19136);
   U916 : BUF_X1 port map( A => n3126, Z => n19137);
   U917 : BUF_X1 port map( A => n3126, Z => n19138);
   U918 : BUF_X1 port map( A => n3009, Z => n19333);
   U919 : BUF_X1 port map( A => n3009, Z => n19334);
   U920 : BUF_X1 port map( A => n3009, Z => n19335);
   U921 : BUF_X1 port map( A => n3009, Z => n19336);
   U922 : BUF_X1 port map( A => n3009, Z => n19337);
   U923 : BUF_X1 port map( A => n3147, Z => n19072);
   U924 : BUF_X1 port map( A => n3147, Z => n19068);
   U925 : BUF_X1 port map( A => n3147, Z => n19069);
   U926 : BUF_X1 port map( A => n3147, Z => n19070);
   U927 : BUF_X1 port map( A => n3147, Z => n19071);
   U928 : BUF_X1 port map( A => n3010, Z => n19327);
   U929 : BUF_X1 port map( A => n3010, Z => n19328);
   U930 : BUF_X1 port map( A => n3010, Z => n19329);
   U931 : BUF_X1 port map( A => n3010, Z => n19330);
   U932 : BUF_X1 port map( A => n3010, Z => n19331);
   U933 : BUF_X1 port map( A => n3127, Z => n19128);
   U934 : BUF_X1 port map( A => n3127, Z => n19129);
   U935 : BUF_X1 port map( A => n3127, Z => n19130);
   U936 : BUF_X1 port map( A => n3127, Z => n19131);
   U937 : BUF_X1 port map( A => n3127, Z => n19132);
   U938 : BUF_X1 port map( A => n3159, Z => n19012);
   U939 : BUF_X1 port map( A => n3159, Z => n19008);
   U940 : BUF_X1 port map( A => n3159, Z => n19009);
   U941 : BUF_X1 port map( A => n3159, Z => n19010);
   U942 : BUF_X1 port map( A => n3110, Z => n19201);
   U943 : BUF_X1 port map( A => n3115, Z => n19177);
   U944 : BUF_X1 port map( A => n3105, Z => n19225);
   U945 : BUF_X1 port map( A => n3036, Z => n19249);
   U946 : BUF_X1 port map( A => n2983, Z => n19424);
   U947 : BUF_X1 port map( A => n2990, Z => n19400);
   U948 : BUF_X1 port map( A => n2977, Z => n19448);
   U949 : BUF_X1 port map( A => n2997, Z => n19376);
   U950 : BUF_X1 port map( A => n3110, Z => n19202);
   U951 : BUF_X1 port map( A => n3115, Z => n19178);
   U952 : BUF_X1 port map( A => n3105, Z => n19226);
   U953 : BUF_X1 port map( A => n3036, Z => n19250);
   U954 : BUF_X1 port map( A => n2983, Z => n19425);
   U955 : BUF_X1 port map( A => n2990, Z => n19401);
   U956 : BUF_X1 port map( A => n2977, Z => n19449);
   U957 : BUF_X1 port map( A => n2997, Z => n19377);
   U958 : BUF_X1 port map( A => n3110, Z => n19203);
   U959 : BUF_X1 port map( A => n3115, Z => n19179);
   U960 : BUF_X1 port map( A => n3105, Z => n19227);
   U961 : BUF_X1 port map( A => n3036, Z => n19251);
   U962 : BUF_X1 port map( A => n2983, Z => n19426);
   U963 : BUF_X1 port map( A => n2990, Z => n19402);
   U964 : BUF_X1 port map( A => n2977, Z => n19450);
   U965 : BUF_X1 port map( A => n2997, Z => n19378);
   U966 : BUF_X1 port map( A => n3159, Z => n19011);
   U967 : BUF_X1 port map( A => n3110, Z => n19204);
   U968 : BUF_X1 port map( A => n3115, Z => n19180);
   U969 : BUF_X1 port map( A => n3105, Z => n19228);
   U970 : BUF_X1 port map( A => n3036, Z => n19252);
   U971 : BUF_X1 port map( A => n2983, Z => n19427);
   U972 : BUF_X1 port map( A => n2990, Z => n19403);
   U973 : BUF_X1 port map( A => n2977, Z => n19451);
   U974 : BUF_X1 port map( A => n2997, Z => n19379);
   U975 : BUF_X1 port map( A => n3110, Z => n19205);
   U976 : BUF_X1 port map( A => n3115, Z => n19181);
   U977 : BUF_X1 port map( A => n3105, Z => n19229);
   U978 : BUF_X1 port map( A => n3036, Z => n19253);
   U979 : BUF_X1 port map( A => n2983, Z => n19428);
   U980 : BUF_X1 port map( A => n2990, Z => n19404);
   U981 : BUF_X1 port map( A => n2977, Z => n19452);
   U982 : BUF_X1 port map( A => n2997, Z => n19380);
   U983 : NAND2_X1 port map( A1 => n11635, A2 => n11643, ZN => n3122);
   U984 : NAND2_X1 port map( A1 => n11633, A2 => n11643, ZN => n3112);
   U985 : NAND2_X1 port map( A1 => n11587, A2 => n11601, ZN => n2993);
   U986 : NAND2_X1 port map( A1 => n11589, A2 => n11601, ZN => n3005);
   U987 : BUF_X1 port map( A => n3124, Z => n19146);
   U988 : BUF_X1 port map( A => n3132, Z => n19104);
   U989 : BUF_X1 port map( A => n3137, Z => n19080);
   U990 : BUF_X1 port map( A => n3124, Z => n19147);
   U991 : BUF_X1 port map( A => n3132, Z => n19105);
   U992 : BUF_X1 port map( A => n3137, Z => n19081);
   U993 : BUF_X1 port map( A => n3124, Z => n19148);
   U994 : BUF_X1 port map( A => n3132, Z => n19106);
   U995 : BUF_X1 port map( A => n3137, Z => n19082);
   U996 : BUF_X1 port map( A => n3124, Z => n19149);
   U997 : BUF_X1 port map( A => n3132, Z => n19107);
   U998 : BUF_X1 port map( A => n3137, Z => n19083);
   U999 : BUF_X1 port map( A => n3124, Z => n19150);
   U1000 : BUF_X1 port map( A => n3132, Z => n19108);
   U1001 : BUF_X1 port map( A => n3137, Z => n19084);
   U1002 : BUF_X1 port map( A => n3120, Z => n19171);
   U1003 : BUF_X1 port map( A => n3015, Z => n19303);
   U1004 : BUF_X1 port map( A => n3007, Z => n19345);
   U1005 : BUF_X1 port map( A => n3003, Z => n19370);
   U1006 : BUF_X1 port map( A => n3022, Z => n19279);
   U1007 : BUF_X1 port map( A => n3120, Z => n19172);
   U1008 : BUF_X1 port map( A => n3015, Z => n19304);
   U1009 : BUF_X1 port map( A => n3007, Z => n19346);
   U1010 : BUF_X1 port map( A => n3003, Z => n19371);
   U1011 : BUF_X1 port map( A => n3022, Z => n19280);
   U1012 : BUF_X1 port map( A => n3120, Z => n19173);
   U1013 : BUF_X1 port map( A => n3015, Z => n19305);
   U1014 : BUF_X1 port map( A => n3007, Z => n19347);
   U1015 : BUF_X1 port map( A => n3003, Z => n19372);
   U1016 : BUF_X1 port map( A => n3022, Z => n19281);
   U1017 : BUF_X1 port map( A => n3120, Z => n19174);
   U1018 : BUF_X1 port map( A => n3015, Z => n19306);
   U1019 : BUF_X1 port map( A => n3007, Z => n19348);
   U1020 : BUF_X1 port map( A => n3003, Z => n19373);
   U1021 : BUF_X1 port map( A => n3022, Z => n19282);
   U1022 : BUF_X1 port map( A => n3120, Z => n19175);
   U1023 : BUF_X1 port map( A => n3015, Z => n19307);
   U1024 : BUF_X1 port map( A => n3007, Z => n19349);
   U1025 : BUF_X1 port map( A => n3003, Z => n19374);
   U1026 : BUF_X1 port map( A => n3022, Z => n19283);
   U1027 : BUF_X1 port map( A => n3198, Z => n18922);
   U1028 : BUF_X1 port map( A => n3198, Z => n18918);
   U1029 : BUF_X1 port map( A => n3198, Z => n18919);
   U1030 : BUF_X1 port map( A => n3198, Z => n18920);
   U1031 : BUF_X1 port map( A => n3198, Z => n18921);
   U1032 : BUF_X1 port map( A => n3123, Z => n19152);
   U1033 : BUF_X1 port map( A => n3008, Z => n19339);
   U1034 : BUF_X1 port map( A => n3006, Z => n19351);
   U1035 : BUF_X1 port map( A => n3123, Z => n19153);
   U1036 : BUF_X1 port map( A => n3008, Z => n19340);
   U1037 : BUF_X1 port map( A => n3006, Z => n19352);
   U1038 : BUF_X1 port map( A => n3123, Z => n19154);
   U1039 : BUF_X1 port map( A => n3008, Z => n19341);
   U1040 : BUF_X1 port map( A => n3006, Z => n19353);
   U1041 : BUF_X1 port map( A => n3123, Z => n19155);
   U1042 : BUF_X1 port map( A => n3008, Z => n19342);
   U1043 : BUF_X1 port map( A => n3006, Z => n19354);
   U1044 : BUF_X1 port map( A => n3123, Z => n19156);
   U1045 : BUF_X1 port map( A => n3008, Z => n19343);
   U1046 : BUF_X1 port map( A => n3006, Z => n19355);
   U1047 : BUF_X1 port map( A => n3125, Z => n19140);
   U1048 : BUF_X1 port map( A => n3133, Z => n19098);
   U1049 : BUF_X1 port map( A => n3138, Z => n19074);
   U1050 : BUF_X1 port map( A => n3016, Z => n19297);
   U1051 : BUF_X1 port map( A => n3023, Z => n19273);
   U1052 : BUF_X1 port map( A => n3125, Z => n19141);
   U1053 : BUF_X1 port map( A => n3133, Z => n19099);
   U1054 : BUF_X1 port map( A => n3138, Z => n19075);
   U1055 : BUF_X1 port map( A => n3016, Z => n19298);
   U1056 : BUF_X1 port map( A => n3023, Z => n19274);
   U1057 : BUF_X1 port map( A => n3125, Z => n19142);
   U1058 : BUF_X1 port map( A => n3133, Z => n19100);
   U1059 : BUF_X1 port map( A => n3138, Z => n19076);
   U1060 : BUF_X1 port map( A => n3016, Z => n19299);
   U1061 : BUF_X1 port map( A => n3023, Z => n19275);
   U1062 : BUF_X1 port map( A => n3125, Z => n19143);
   U1063 : BUF_X1 port map( A => n3133, Z => n19101);
   U1064 : BUF_X1 port map( A => n3138, Z => n19077);
   U1065 : BUF_X1 port map( A => n3016, Z => n19300);
   U1066 : BUF_X1 port map( A => n3023, Z => n19276);
   U1067 : BUF_X1 port map( A => n3125, Z => n19144);
   U1068 : BUF_X1 port map( A => n3133, Z => n19102);
   U1069 : BUF_X1 port map( A => n3138, Z => n19078);
   U1070 : BUF_X1 port map( A => n3016, Z => n19301);
   U1071 : BUF_X1 port map( A => n3023, Z => n19277);
   U1072 : BUF_X1 port map( A => n3107, Z => n19213);
   U1073 : BUF_X1 port map( A => n3107, Z => n19214);
   U1074 : BUF_X1 port map( A => n3107, Z => n19215);
   U1075 : BUF_X1 port map( A => n3107, Z => n19216);
   U1076 : BUF_X1 port map( A => n3107, Z => n19217);
   U1077 : BUF_X1 port map( A => n3102, Z => n19237);
   U1078 : BUF_X1 port map( A => n2980, Z => n19436);
   U1079 : BUF_X1 port map( A => n2986, Z => n19412);
   U1080 : BUF_X1 port map( A => n3102, Z => n19238);
   U1081 : BUF_X1 port map( A => n2980, Z => n19437);
   U1082 : BUF_X1 port map( A => n2986, Z => n19413);
   U1083 : BUF_X1 port map( A => n3102, Z => n19239);
   U1084 : BUF_X1 port map( A => n2980, Z => n19438);
   U1085 : BUF_X1 port map( A => n2986, Z => n19414);
   U1086 : BUF_X1 port map( A => n3102, Z => n19240);
   U1087 : BUF_X1 port map( A => n2980, Z => n19439);
   U1088 : BUF_X1 port map( A => n2986, Z => n19415);
   U1089 : BUF_X1 port map( A => n3102, Z => n19241);
   U1090 : BUF_X1 port map( A => n2980, Z => n19440);
   U1091 : BUF_X1 port map( A => n2986, Z => n19416);
   U1092 : BUF_X1 port map( A => n3161, Z => n19000);
   U1093 : BUF_X1 port map( A => n3156, Z => n19024);
   U1094 : BUF_X1 port map( A => n3161, Z => n18996);
   U1095 : BUF_X1 port map( A => n3156, Z => n19020);
   U1096 : BUF_X1 port map( A => n3161, Z => n18997);
   U1097 : BUF_X1 port map( A => n3156, Z => n19021);
   U1098 : BUF_X1 port map( A => n3161, Z => n18998);
   U1099 : BUF_X1 port map( A => n3156, Z => n19022);
   U1100 : BUF_X1 port map( A => n3161, Z => n18999);
   U1101 : BUF_X1 port map( A => n3156, Z => n19023);
   U1102 : BUF_X1 port map( A => n3106, Z => n19219);
   U1103 : BUF_X1 port map( A => n2985, Z => n19418);
   U1104 : BUF_X1 port map( A => n2780, Z => n19466);
   U1105 : BUF_X1 port map( A => n3032, Z => n19267);
   U1106 : BUF_X1 port map( A => n3111, Z => n19195);
   U1107 : BUF_X1 port map( A => n3037, Z => n19243);
   U1108 : BUF_X1 port map( A => n2979, Z => n19442);
   U1109 : BUF_X1 port map( A => n2992, Z => n19394);
   U1110 : AND2_X1 port map( A1 => n11652, A2 => n11643, ZN => n3135);
   U1111 : AND2_X1 port map( A1 => n11643, A2 => n11642, ZN => n3114);
   U1112 : AND2_X1 port map( A1 => n11611, A2 => n11601, ZN => n3019);
   U1113 : AND2_X1 port map( A1 => n11601, A2 => n11600, ZN => n2995);
   U1114 : AND2_X1 port map( A1 => n11682, A2 => n11681, ZN => n11670);
   U1115 : INV_X1 port map( A => n11686, ZN => n11677);
   U1116 : BUF_X1 port map( A => n3004, Z => n19363);
   U1117 : BUF_X1 port map( A => n3121, Z => n19164);
   U1118 : BUF_X1 port map( A => n3004, Z => n19364);
   U1119 : BUF_X1 port map( A => n3121, Z => n19165);
   U1120 : BUF_X1 port map( A => n1873, Z => n19994);
   U1121 : BUF_X1 port map( A => n1873, Z => n19995);
   U1122 : BUF_X1 port map( A => n1945, Z => n19938);
   U1123 : BUF_X1 port map( A => n1945, Z => n19939);
   U1124 : BUF_X1 port map( A => n2017, Z => n19882);
   U1125 : BUF_X1 port map( A => n2017, Z => n19883);
   U1126 : BUF_X1 port map( A => n2243, Z => n19658);
   U1127 : BUF_X1 port map( A => n2243, Z => n19659);
   U1128 : BUF_X1 port map( A => n2198, Z => n19770);
   U1129 : BUF_X1 port map( A => n2198, Z => n19771);
   U1130 : BUF_X1 port map( A => n2443, Z => n19546);
   U1131 : BUF_X1 port map( A => n2443, Z => n19547);
   U1132 : BUF_X1 port map( A => n1729, Z => n20106);
   U1133 : BUF_X1 port map( A => n1703, Z => n20330);
   U1134 : BUF_X1 port map( A => n1718, Z => n20218);
   U1135 : BUF_X1 port map( A => n1729, Z => n20107);
   U1136 : BUF_X1 port map( A => n1703, Z => n20331);
   U1137 : BUF_X1 port map( A => n1718, Z => n20219);
   U1138 : BUF_X1 port map( A => n1865, Z => n20050);
   U1139 : BUF_X1 port map( A => n1723, Z => n20162);
   U1140 : BUF_X1 port map( A => n1865, Z => n20051);
   U1141 : BUF_X1 port map( A => n1723, Z => n20163);
   U1142 : BUF_X1 port map( A => n1711, Z => n20274);
   U1143 : BUF_X1 port map( A => n1711, Z => n20275);
   U1144 : BUF_X1 port map( A => n2089, Z => n19826);
   U1145 : BUF_X1 port map( A => n2089, Z => n19827);
   U1146 : BUF_X1 port map( A => n2258, Z => n19602);
   U1147 : BUF_X1 port map( A => n2258, Z => n19603);
   U1148 : BUF_X1 port map( A => n2213, Z => n19714);
   U1149 : BUF_X1 port map( A => n2213, Z => n19715);
   U1150 : BUF_X1 port map( A => n19966, Z => n19964);
   U1151 : BUF_X1 port map( A => n19966, Z => n19963);
   U1152 : BUF_X1 port map( A => n19967, Z => n19962);
   U1153 : BUF_X1 port map( A => n19967, Z => n19961);
   U1154 : BUF_X1 port map( A => n19967, Z => n19960);
   U1155 : BUF_X1 port map( A => n20022, Z => n20020);
   U1156 : BUF_X1 port map( A => n20022, Z => n20019);
   U1157 : BUF_X1 port map( A => n20023, Z => n20018);
   U1158 : BUF_X1 port map( A => n20023, Z => n20017);
   U1159 : BUF_X1 port map( A => n20023, Z => n20016);
   U1160 : BUF_X1 port map( A => n19798, Z => n19796);
   U1161 : BUF_X1 port map( A => n19798, Z => n19795);
   U1162 : BUF_X1 port map( A => n19799, Z => n19794);
   U1163 : BUF_X1 port map( A => n19799, Z => n19793);
   U1164 : BUF_X1 port map( A => n19799, Z => n19792);
   U1165 : BUF_X1 port map( A => n19686, Z => n19684);
   U1166 : BUF_X1 port map( A => n19686, Z => n19683);
   U1167 : BUF_X1 port map( A => n19687, Z => n19682);
   U1168 : BUF_X1 port map( A => n19687, Z => n19681);
   U1169 : BUF_X1 port map( A => n19687, Z => n19680);
   U1170 : BUF_X1 port map( A => n19910, Z => n19908);
   U1171 : BUF_X1 port map( A => n19910, Z => n19907);
   U1172 : BUF_X1 port map( A => n19911, Z => n19906);
   U1173 : BUF_X1 port map( A => n19911, Z => n19905);
   U1174 : BUF_X1 port map( A => n19911, Z => n19904);
   U1175 : BUF_X1 port map( A => n19630, Z => n19628);
   U1176 : BUF_X1 port map( A => n19630, Z => n19627);
   U1177 : BUF_X1 port map( A => n19631, Z => n19626);
   U1178 : BUF_X1 port map( A => n19631, Z => n19625);
   U1179 : BUF_X1 port map( A => n19631, Z => n19624);
   U1180 : BUF_X1 port map( A => n19854, Z => n19852);
   U1181 : BUF_X1 port map( A => n19854, Z => n19851);
   U1182 : BUF_X1 port map( A => n19855, Z => n19850);
   U1183 : BUF_X1 port map( A => n19855, Z => n19849);
   U1184 : BUF_X1 port map( A => n19855, Z => n19848);
   U1185 : BUF_X1 port map( A => n19742, Z => n19740);
   U1186 : BUF_X1 port map( A => n19742, Z => n19739);
   U1187 : BUF_X1 port map( A => n19743, Z => n19738);
   U1188 : BUF_X1 port map( A => n19743, Z => n19737);
   U1189 : BUF_X1 port map( A => n19743, Z => n19736);
   U1190 : BUF_X1 port map( A => n20134, Z => n20132);
   U1191 : BUF_X1 port map( A => n20134, Z => n20131);
   U1192 : BUF_X1 port map( A => n20135, Z => n20130);
   U1193 : BUF_X1 port map( A => n20135, Z => n20129);
   U1194 : BUF_X1 port map( A => n20135, Z => n20128);
   U1195 : BUF_X1 port map( A => n20078, Z => n20076);
   U1196 : BUF_X1 port map( A => n20078, Z => n20075);
   U1197 : BUF_X1 port map( A => n20079, Z => n20074);
   U1198 : BUF_X1 port map( A => n20079, Z => n20073);
   U1199 : BUF_X1 port map( A => n20079, Z => n20072);
   U1200 : BUF_X1 port map( A => n20302, Z => n20300);
   U1201 : BUF_X1 port map( A => n20302, Z => n20299);
   U1202 : BUF_X1 port map( A => n20303, Z => n20298);
   U1203 : BUF_X1 port map( A => n20303, Z => n20297);
   U1204 : BUF_X1 port map( A => n20303, Z => n20296);
   U1205 : BUF_X1 port map( A => n20190, Z => n20188);
   U1206 : BUF_X1 port map( A => n20190, Z => n20187);
   U1207 : BUF_X1 port map( A => n20191, Z => n20186);
   U1208 : BUF_X1 port map( A => n20191, Z => n20185);
   U1209 : BUF_X1 port map( A => n20191, Z => n20184);
   U1210 : BUF_X1 port map( A => n20550, Z => n20548);
   U1211 : BUF_X1 port map( A => n20550, Z => n20547);
   U1212 : BUF_X1 port map( A => n20551, Z => n20546);
   U1213 : BUF_X1 port map( A => n20551, Z => n20545);
   U1214 : BUF_X1 port map( A => n20551, Z => n20544);
   U1215 : BUF_X1 port map( A => n20246, Z => n20244);
   U1216 : BUF_X1 port map( A => n20246, Z => n20243);
   U1217 : BUF_X1 port map( A => n20247, Z => n20242);
   U1218 : BUF_X1 port map( A => n20247, Z => n20241);
   U1219 : BUF_X1 port map( A => n20247, Z => n20240);
   U1220 : BUF_X1 port map( A => n19574, Z => n19572);
   U1221 : BUF_X1 port map( A => n19574, Z => n19571);
   U1222 : BUF_X1 port map( A => n19575, Z => n19570);
   U1223 : BUF_X1 port map( A => n19575, Z => n19569);
   U1224 : BUF_X1 port map( A => n19575, Z => n19568);
   U1225 : BUF_X1 port map( A => n19518, Z => n19516);
   U1226 : BUF_X1 port map( A => n19518, Z => n19515);
   U1227 : BUF_X1 port map( A => n19519, Z => n19514);
   U1228 : BUF_X1 port map( A => n19519, Z => n19513);
   U1229 : BUF_X1 port map( A => n19519, Z => n19512);
   U1230 : BUF_X1 port map( A => n2767, Z => n19490);
   U1231 : BUF_X1 port map( A => n2767, Z => n19491);
   U1232 : BUF_X1 port map( A => n19966, Z => n19965);
   U1233 : BUF_X1 port map( A => n20022, Z => n20021);
   U1234 : BUF_X1 port map( A => n19798, Z => n19797);
   U1235 : BUF_X1 port map( A => n19686, Z => n19685);
   U1236 : BUF_X1 port map( A => n19910, Z => n19909);
   U1237 : BUF_X1 port map( A => n19630, Z => n19629);
   U1238 : BUF_X1 port map( A => n19742, Z => n19741);
   U1239 : BUF_X1 port map( A => n19854, Z => n19853);
   U1240 : BUF_X1 port map( A => n20134, Z => n20133);
   U1241 : BUF_X1 port map( A => n20078, Z => n20077);
   U1242 : BUF_X1 port map( A => n20302, Z => n20301);
   U1243 : BUF_X1 port map( A => n20190, Z => n20189);
   U1244 : BUF_X1 port map( A => n20550, Z => n20549);
   U1245 : BUF_X1 port map( A => n20246, Z => n20245);
   U1246 : BUF_X1 port map( A => n19574, Z => n19573);
   U1247 : BUF_X1 port map( A => n19518, Z => n19517);
   U1248 : OAI211_X1 port map( C1 => n2216, C2 => n11681, A => n11682, B => 
                           n11715, ZN => n3198);
   U1249 : NOR3_X1 port map( A1 => n11653, A2 => n11654, A3 => n11655, ZN => 
                           n11635);
   U1250 : NOR3_X1 port map( A1 => n11563, A2 => n11653, A3 => n11655, ZN => 
                           n11633);
   U1251 : NOR3_X1 port map( A1 => n11614, A2 => n11612, A3 => n11613, ZN => 
                           n11587);
   U1252 : NOR3_X1 port map( A1 => n11574, A2 => n11612, A3 => n11613, ZN => 
                           n11589);
   U1253 : BUF_X1 port map( A => n3170, Z => n18973);
   U1254 : BUF_X1 port map( A => n3170, Z => n18974);
   U1255 : NOR3_X1 port map( A1 => n11614, A2 => n11573, A3 => n11613, ZN => 
                           n11600);
   U1256 : BUF_X1 port map( A => n3172, Z => n18967);
   U1257 : BUF_X1 port map( A => n3172, Z => n18968);
   U1258 : BUF_X1 port map( A => n3172, Z => n18969);
   U1259 : NOR3_X1 port map( A1 => n11573, A2 => n11574, A3 => n11613, ZN => 
                           n11611);
   U1260 : BUF_X1 port map( A => n3174, Z => n18964);
   U1261 : BUF_X1 port map( A => n3174, Z => n18960);
   U1262 : BUF_X1 port map( A => n3174, Z => n18961);
   U1263 : BUF_X1 port map( A => n3174, Z => n18962);
   U1264 : BUF_X1 port map( A => n3174, Z => n18963);
   U1265 : BUF_X1 port map( A => n3149, Z => n19060);
   U1266 : BUF_X1 port map( A => n3149, Z => n19056);
   U1267 : BUF_X1 port map( A => n3149, Z => n19057);
   U1268 : BUF_X1 port map( A => n3149, Z => n19058);
   U1269 : BUF_X1 port map( A => n3149, Z => n19059);
   U1270 : BUF_X1 port map( A => n3148, Z => n19066);
   U1271 : BUF_X1 port map( A => n3148, Z => n19062);
   U1272 : BUF_X1 port map( A => n3148, Z => n19063);
   U1273 : BUF_X1 port map( A => n3148, Z => n19064);
   U1274 : BUF_X1 port map( A => n3148, Z => n19065);
   U1275 : NOR3_X1 port map( A1 => n18915, A2 => n11716, A3 => n11674, ZN => 
                           n11682);
   U1276 : NAND2_X1 port map( A1 => n11644, A2 => n11634, ZN => n3124);
   U1277 : NAND2_X1 port map( A1 => n11645, A2 => n11643, ZN => n3107);
   U1278 : NAND2_X1 port map( A1 => n11645, A2 => n11634, ZN => n3132);
   U1279 : NAND2_X1 port map( A1 => n11645, A2 => n11636, ZN => n3137);
   U1280 : OAI221_X1 port map( B1 => n1699, B2 => n1797, C1 => n1705, C2 => 
                           n1726, A => n20352, ZN => n1729);
   U1281 : OAI221_X1 port map( B1 => n1699, B2 => n1704, C1 => n1698, C2 => 
                           n1705, A => n20352, ZN => n1703);
   U1282 : OAI221_X1 port map( B1 => n1699, B2 => n1719, C1 => n1705, C2 => 
                           n1715, A => n20352, ZN => n1718);
   U1283 : OAI221_X1 port map( B1 => n1709, B2 => n1797, C1 => n1712, C2 => 
                           n1726, A => n20352, ZN => n1865);
   U1284 : OAI221_X1 port map( B1 => n1709, B2 => n1719, C1 => n1712, C2 => 
                           n1715, A => n20353, ZN => n1723);
   U1285 : OAI221_X1 port map( B1 => n1704, B2 => n1709, C1 => n1698, C2 => 
                           n1712, A => n20352, ZN => n1711);
   U1286 : OAI221_X1 port map( B1 => n1704, B2 => n2085, C1 => n1698, C2 => 
                           n2090, A => n20353, ZN => n2089);
   U1287 : OAI221_X1 port map( B1 => n1797, B2 => n2085, C1 => n1726, C2 => 
                           n2090, A => n20354, ZN => n2258);
   U1288 : NAND2_X1 port map( A1 => n11642, A2 => n11634, ZN => n3123);
   U1289 : NAND2_X1 port map( A1 => n11652, A2 => n11634, ZN => n3120);
   U1290 : NAND2_X1 port map( A1 => n11652, A2 => n11636, ZN => n3138);
   U1291 : OAI221_X1 port map( B1 => n1719, B2 => n2085, C1 => n1715, C2 => 
                           n2090, A => n20353, ZN => n2213);
   U1292 : BUF_X1 port map( A => n3153, Z => n19042);
   U1293 : BUF_X1 port map( A => n3153, Z => n19038);
   U1294 : BUF_X1 port map( A => n3153, Z => n19039);
   U1295 : BUF_X1 port map( A => n3153, Z => n19040);
   U1296 : BUF_X1 port map( A => n3153, Z => n19041);
   U1297 : BUF_X1 port map( A => n3163, Z => n18994);
   U1298 : BUF_X1 port map( A => n3180, Z => n18952);
   U1299 : BUF_X1 port map( A => n3163, Z => n18990);
   U1300 : BUF_X1 port map( A => n3180, Z => n18948);
   U1301 : BUF_X1 port map( A => n3163, Z => n18991);
   U1302 : BUF_X1 port map( A => n3180, Z => n18949);
   U1303 : BUF_X1 port map( A => n3163, Z => n18992);
   U1304 : BUF_X1 port map( A => n3180, Z => n18950);
   U1305 : BUF_X1 port map( A => n3163, Z => n18993);
   U1306 : BUF_X1 port map( A => n3180, Z => n18951);
   U1307 : BUF_X1 port map( A => n3190, Z => n18934);
   U1308 : BUF_X1 port map( A => n3190, Z => n18930);
   U1309 : BUF_X1 port map( A => n3190, Z => n18931);
   U1310 : BUF_X1 port map( A => n3190, Z => n18932);
   U1311 : BUF_X1 port map( A => n3190, Z => n18933);
   U1312 : BUF_X1 port map( A => n3150, Z => n19054);
   U1313 : BUF_X1 port map( A => n3155, Z => n19030);
   U1314 : BUF_X1 port map( A => n3150, Z => n19051);
   U1315 : BUF_X1 port map( A => n3155, Z => n19027);
   U1316 : BUF_X1 port map( A => n3150, Z => n19052);
   U1317 : BUF_X1 port map( A => n3155, Z => n19028);
   U1318 : BUF_X1 port map( A => n3155, Z => n19029);
   U1319 : NAND2_X1 port map( A1 => n1947, A2 => n2764, ZN => n2085);
   U1320 : BUF_X1 port map( A => n3202, Z => n18913);
   U1321 : BUF_X1 port map( A => n3202, Z => n18910);
   U1322 : BUF_X1 port map( A => n3202, Z => n18911);
   U1323 : BUF_X1 port map( A => n3202, Z => n18912);
   U1324 : BUF_X1 port map( A => n3150, Z => n19053);
   U1325 : BUF_X1 port map( A => n3176, Z => n18958);
   U1326 : BUF_X1 port map( A => n3176, Z => n18954);
   U1327 : BUF_X1 port map( A => n3176, Z => n18955);
   U1328 : BUF_X1 port map( A => n3176, Z => n18956);
   U1329 : BUF_X1 port map( A => n3176, Z => n18957);
   U1330 : BUF_X1 port map( A => n3154, Z => n19036);
   U1331 : BUF_X1 port map( A => n3165, Z => n18988);
   U1332 : BUF_X1 port map( A => n3184, Z => n18946);
   U1333 : BUF_X1 port map( A => n3154, Z => n19032);
   U1334 : BUF_X1 port map( A => n3165, Z => n18984);
   U1335 : BUF_X1 port map( A => n3184, Z => n18942);
   U1336 : BUF_X1 port map( A => n3154, Z => n19033);
   U1337 : BUF_X1 port map( A => n3165, Z => n18985);
   U1338 : BUF_X1 port map( A => n3184, Z => n18943);
   U1339 : BUF_X1 port map( A => n3154, Z => n19034);
   U1340 : BUF_X1 port map( A => n3165, Z => n18986);
   U1341 : BUF_X1 port map( A => n3184, Z => n18944);
   U1342 : BUF_X1 port map( A => n3154, Z => n19035);
   U1343 : BUF_X1 port map( A => n3165, Z => n18987);
   U1344 : BUF_X1 port map( A => n3184, Z => n18945);
   U1345 : NOR2_X1 port map( A1 => n11736, A2 => n11702, ZN => n11724);
   U1346 : AND3_X1 port map( A1 => n11660, A2 => n11565, A3 => n11658, ZN => 
                           n11643);
   U1347 : AND3_X1 port map( A1 => n11621, A2 => n11616, A3 => n11617, ZN => 
                           n11601);
   U1348 : BUF_X1 port map( A => n3172, Z => n18966);
   U1349 : NAND2_X1 port map( A1 => n11602, A2 => n11588, ZN => n3007);
   U1350 : BUF_X1 port map( A => n3166, Z => n18982);
   U1351 : BUF_X1 port map( A => n3166, Z => n18978);
   U1352 : BUF_X1 port map( A => n3166, Z => n18979);
   U1353 : BUF_X1 port map( A => n3166, Z => n18980);
   U1354 : BUF_X1 port map( A => n3166, Z => n18981);
   U1355 : BUF_X1 port map( A => n3160, Z => n19006);
   U1356 : BUF_X1 port map( A => n3160, Z => n19002);
   U1357 : BUF_X1 port map( A => n3160, Z => n19003);
   U1358 : BUF_X1 port map( A => n3160, Z => n19004);
   U1359 : BUF_X1 port map( A => n3160, Z => n19005);
   U1360 : NAND2_X1 port map( A1 => n11603, A2 => n11601, ZN => n2986);
   U1361 : NAND2_X1 port map( A1 => n11603, A2 => n11588, ZN => n3015);
   U1362 : NAND2_X1 port map( A1 => n11603, A2 => n11590, ZN => n3022);
   U1363 : NAND2_X1 port map( A1 => n11635, A2 => n11634, ZN => n3102);
   U1364 : NAND2_X1 port map( A1 => n11633, A2 => n11639, ZN => n3133);
   U1365 : NAND2_X1 port map( A1 => n11589, A2 => n11588, ZN => n2980);
   U1366 : NAND2_X1 port map( A1 => n11587, A2 => n11594, ZN => n3016);
   U1367 : BUF_X1 port map( A => n3170, Z => n18976);
   U1368 : BUF_X1 port map( A => n3170, Z => n18975);
   U1369 : BUF_X1 port map( A => n3196, Z => n18928);
   U1370 : BUF_X1 port map( A => n3196, Z => n18924);
   U1371 : BUF_X1 port map( A => n3196, Z => n18925);
   U1372 : BUF_X1 port map( A => n3196, Z => n18926);
   U1373 : BUF_X1 port map( A => n3196, Z => n18927);
   U1374 : NAND2_X1 port map( A1 => n11642, A2 => n11636, ZN => n3128);
   U1375 : BUF_X1 port map( A => n3206, Z => n18907);
   U1376 : BUF_X1 port map( A => n3206, Z => n18903);
   U1377 : BUF_X1 port map( A => n3206, Z => n18904);
   U1378 : BUF_X1 port map( A => n3206, Z => n18905);
   U1379 : BUF_X1 port map( A => n3206, Z => n18906);
   U1380 : BUF_X1 port map( A => n3172, Z => n18970);
   U1381 : NAND2_X1 port map( A1 => n11611, A2 => n11588, ZN => n3003);
   U1382 : NAND2_X1 port map( A1 => n11600, A2 => n11588, ZN => n3006);
   U1383 : NAND2_X1 port map( A1 => n11591, A2 => n11594, ZN => n3008);
   U1384 : NAND2_X1 port map( A1 => n11637, A2 => n11639, ZN => n3125);
   U1385 : NOR2_X1 port map( A1 => n18917, A2 => n2090, ZN => n11711);
   U1386 : NAND2_X1 port map( A1 => n11611, A2 => n11590, ZN => n3023);
   U1387 : NAND2_X1 port map( A1 => n11692, A2 => n11679, ZN => n3161);
   U1388 : NAND2_X1 port map( A1 => n11676, A2 => n11679, ZN => n3156);
   U1389 : BUF_X1 port map( A => n3151, Z => n19048);
   U1390 : BUF_X1 port map( A => n3151, Z => n19044);
   U1391 : BUF_X1 port map( A => n3151, Z => n19045);
   U1392 : BUF_X1 port map( A => n3151, Z => n19046);
   U1393 : BUF_X2 port map( A => n3151, Z => n19047);
   U1394 : BUF_X1 port map( A => n3150, Z => n19050);
   U1395 : BUF_X1 port map( A => n3155, Z => n19026);
   U1396 : NOR2_X1 port map( A1 => n18916, A2 => n11702, ZN => n11718);
   U1397 : INV_X1 port map( A => n11671, ZN => n11688);
   U1398 : BUF_X1 port map( A => n3202, Z => n18909);
   U1399 : NAND2_X1 port map( A1 => n11639, A2 => n11644, ZN => n3106);
   U1400 : INV_X1 port map( A => n11708, ZN => n11679);
   U1401 : NAND2_X1 port map( A1 => n11636, A2 => n11644, ZN => n3126);
   U1402 : NAND2_X1 port map( A1 => n11635, A2 => n11639, ZN => n3037);
   U1403 : NAND2_X1 port map( A1 => n11633, A2 => n11636, ZN => n3111);
   U1404 : NAND2_X1 port map( A1 => n11589, A2 => n11594, ZN => n2979);
   U1405 : NAND2_X1 port map( A1 => n11587, A2 => n11590, ZN => n2992);
   U1406 : NAND2_X1 port map( A1 => n11591, A2 => n11588, ZN => n2780);
   U1407 : NAND2_X1 port map( A1 => n11637, A2 => n11634, ZN => n3032);
   U1408 : NAND2_X1 port map( A1 => n11594, A2 => n11602, ZN => n2985);
   U1409 : INV_X1 port map( A => n11574, ZN => n11614);
   U1410 : NAND2_X1 port map( A1 => n11600, A2 => n11590, ZN => n3011);
   U1411 : INV_X1 port map( A => n11573, ZN => n11612);
   U1412 : NAND2_X1 port map( A1 => n11590, A2 => n11602, ZN => n3009);
   U1413 : INV_X1 port map( A => n11654, ZN => n11563);
   U1414 : NAND2_X1 port map( A1 => n11588, A2 => n11596, ZN => n3010);
   U1415 : NAND2_X1 port map( A1 => n11634, A2 => n11640, ZN => n3127);
   U1416 : AND2_X1 port map( A1 => n11645, A2 => n11639, ZN => n3130);
   U1417 : INV_X1 port map( A => n11556, ZN => n2228);
   U1418 : AND2_X1 port map( A1 => n11652, A2 => n11639, ZN => n3129);
   U1419 : AND2_X1 port map( A1 => n11643, A2 => n11644, ZN => n3109);
   U1420 : NAND2_X1 port map( A1 => n11676, A2 => n11677, ZN => n3147);
   U1421 : INV_X1 port map( A => n11710, ZN => n11684);
   U1422 : AND2_X1 port map( A1 => n11639, A2 => n11642, ZN => n3110);
   U1423 : AND2_X1 port map( A1 => n11603, A2 => n11594, ZN => n3013);
   U1424 : AND2_X1 port map( A1 => n11633, A2 => n11634, ZN => n3036);
   U1425 : AND2_X1 port map( A1 => n11635, A2 => n11636, ZN => n3035);
   U1426 : AND2_X1 port map( A1 => n11587, A2 => n11588, ZN => n2977);
   U1427 : AND2_X1 port map( A1 => n11589, A2 => n11590, ZN => n2783);
   U1428 : AND2_X1 port map( A1 => n11591, A2 => n11590, ZN => n2997);
   U1429 : AND2_X1 port map( A1 => n11637, A2 => n11636, ZN => n3115);
   U1430 : AND2_X1 port map( A1 => n11611, A2 => n11594, ZN => n3012);
   U1431 : AND2_X1 port map( A1 => n11601, A2 => n11602, ZN => n2988);
   U1432 : AND2_X1 port map( A1 => n11594, A2 => n11596, ZN => n2983);
   U1433 : AND2_X1 port map( A1 => n11590, A2 => n11596, ZN => n2982);
   U1434 : AND2_X1 port map( A1 => n11639, A2 => n11640, ZN => n3105);
   U1435 : AND2_X1 port map( A1 => n11636, A2 => n11640, ZN => n3104);
   U1436 : AND2_X1 port map( A1 => n11601, A2 => n11591, ZN => n3017);
   U1437 : AND2_X1 port map( A1 => n11594, A2 => n11600, ZN => n2990);
   U1438 : AND2_X1 port map( A1 => n11643, A2 => n11637, ZN => n3134);
   U1439 : AND2_X1 port map( A1 => n11715, A2 => n11684, ZN => n3186);
   U1440 : AND2_X1 port map( A1 => n11676, A2 => n11670, ZN => n3159);
   U1441 : INV_X1 port map( A => n11696, ZN => n11706);
   U1442 : AND2_X1 port map( A1 => n19266, A2 => n20354, ZN => n11658);
   U1443 : AND2_X1 port map( A1 => n19465, A2 => n20354, ZN => n11617);
   U1444 : INV_X1 port map( A => n1946, ZN => n1870);
   U1445 : NAND2_X1 port map( A1 => n11601, A2 => n11596, ZN => n3004);
   U1446 : NAND2_X1 port map( A1 => n11643, A2 => n11640, ZN => n3121);
   U1447 : INV_X1 port map( A => n11692, ZN => n11687);
   U1448 : BUF_X1 port map( A => n1942, Z => n19966);
   U1449 : BUF_X1 port map( A => n1867, Z => n20022);
   U1450 : BUF_X1 port map( A => n1942, Z => n19967);
   U1451 : BUF_X1 port map( A => n1867, Z => n20023);
   U1452 : BUF_X1 port map( A => n2096, Z => n19798);
   U1453 : BUF_X1 port map( A => n2237, Z => n19686);
   U1454 : BUF_X1 port map( A => n2249, Z => n19630);
   U1455 : BUF_X1 port map( A => n2204, Z => n19742);
   U1456 : BUF_X1 port map( A => n2096, Z => n19799);
   U1457 : BUF_X1 port map( A => n2237, Z => n19687);
   U1458 : BUF_X1 port map( A => n2249, Z => n19631);
   U1459 : BUF_X1 port map( A => n2204, Z => n19743);
   U1460 : BUF_X1 port map( A => n1949, Z => n19910);
   U1461 : BUF_X1 port map( A => n2084, Z => n19854);
   U1462 : BUF_X1 port map( A => n1949, Z => n19911);
   U1463 : BUF_X1 port map( A => n2084, Z => n19855);
   U1464 : BUF_X1 port map( A => n1725, Z => n20134);
   U1465 : BUF_X1 port map( A => n1633, Z => n20550);
   U1466 : BUF_X1 port map( A => n1714, Z => n20246);
   U1467 : BUF_X1 port map( A => n1725, Z => n20135);
   U1468 : BUF_X1 port map( A => n1633, Z => n20551);
   U1469 : BUF_X1 port map( A => n1714, Z => n20247);
   U1470 : BUF_X1 port map( A => n1799, Z => n20078);
   U1471 : BUF_X1 port map( A => n1721, Z => n20190);
   U1472 : BUF_X1 port map( A => n1799, Z => n20079);
   U1473 : BUF_X1 port map( A => n1721, Z => n20191);
   U1474 : BUF_X1 port map( A => n1707, Z => n20302);
   U1475 : BUF_X1 port map( A => n1707, Z => n20303);
   U1476 : BUF_X1 port map( A => n2377, Z => n19574);
   U1477 : BUF_X1 port map( A => n2766, Z => n19518);
   U1478 : BUF_X1 port map( A => n2377, Z => n19575);
   U1479 : BUF_X1 port map( A => n2766, Z => n19519);
   U1480 : OAI221_X1 port map( B1 => n1938, B2 => n2085, C1 => n1868, C2 => 
                           n2090, A => n20354, ZN => n2767);
   U1481 : BUF_X1 port map( A => n2781, Z => n19464);
   U1482 : BUF_X1 port map( A => n2781, Z => n19463);
   U1483 : BUF_X1 port map( A => n2781, Z => n19462);
   U1484 : BUF_X1 port map( A => n2781, Z => n19461);
   U1485 : BUF_X1 port map( A => n2781, Z => n19460);
   U1486 : INV_X1 port map( A => n11711, ZN => n11709);
   U1487 : OAI22_X1 port map( A1 => n2015, A2 => n11694, B1 => n11708, B2 => 
                           n11699, ZN => n3206);
   U1488 : AOI21_X1 port map( B1 => n11622, B2 => sub_105_carry_4_port, A => 
                           n11623, ZN => n11574);
   U1489 : OAI21_X1 port map( B1 => U3_U4_Z_0, B2 => n11623, A => 
                           sub_105_carry_4_port, ZN => n11573);
   U1490 : NOR3_X1 port map( A1 => n11573, A2 => N113, A3 => n11614, ZN => 
                           n11602);
   U1491 : OAI211_X1 port map( C1 => n2091, C2 => n11681, A => n11682, B => 
                           n11683, ZN => n3151);
   U1492 : NOR3_X1 port map( A1 => n11574, A2 => N113, A3 => n11573, ZN => 
                           n11603);
   U1493 : NOR3_X1 port map( A1 => n11612, A2 => N113, A3 => n11574, ZN => 
                           n11596);
   U1494 : NOR3_X1 port map( A1 => n11654, A2 => N78, A3 => n11653, ZN => 
                           n11640);
   U1495 : NOR3_X1 port map( A1 => n11612, A2 => N113, A3 => n11614, ZN => 
                           n11591);
   U1496 : NOR3_X1 port map( A1 => n11653, A2 => N78, A3 => n11563, ZN => 
                           n11637);
   U1497 : OAI22_X1 port map( A1 => n11724, A2 => n11723, B1 => n11727, B2 => 
                           n11728, ZN => n11725);
   U1498 : NOR2_X1 port map( A1 => n11729, A2 => n11730, ZN => n11727);
   U1499 : INV_X1 port map( A => n11724, ZN => n11730);
   U1500 : NAND4_X1 port map( A1 => n11670, A2 => n11671, A3 => n11672, A4 => 
                           n1939, ZN => n3149);
   U1501 : NAND4_X1 port map( A1 => n11679, A2 => n11671, A3 => n11672, A4 => 
                           n1939, ZN => n3174);
   U1502 : NOR3_X1 port map( A1 => n1939, A2 => n11688, A3 => n11672, ZN => 
                           n11692);
   U1503 : OAI21_X1 port map( B1 => n11686, B2 => n11699, A => n11721, ZN => 
                           n3202);
   U1504 : OR3_X1 port map( A1 => n2015, A2 => n2375, A3 => n18917, ZN => 
                           n11721);
   U1505 : OAI221_X1 port map( B1 => n1716, B2 => n2014, C1 => n1715, C2 => 
                           n2015, A => n20353, ZN => n2096);
   U1506 : OAI221_X1 port map( B1 => n1727, B2 => n2014, C1 => n1726, C2 => 
                           n2015, A => n20354, ZN => n2237);
   U1507 : OAI221_X1 port map( B1 => n1727, B2 => n2085, C1 => n1726, C2 => 
                           n2086, A => n20354, ZN => n2249);
   U1508 : OAI221_X1 port map( B1 => n1716, B2 => n2085, C1 => n1715, C2 => 
                           n2086, A => n20353, ZN => n2204);
   U1509 : NOR2_X1 port map( A1 => n11726, A2 => n11559, ZN => n11702);
   U1510 : OAI221_X1 port map( B1 => n1700, B2 => n2014, C1 => n1698, C2 => 
                           n2015, A => n20353, ZN => n1949);
   U1511 : OAI221_X1 port map( B1 => n1700, B2 => n2085, C1 => n1698, C2 => 
                           n2086, A => n20353, ZN => n2084);
   U1512 : INV_X1 port map( A => n11707, ZN => n3176);
   U1513 : OAI21_X1 port map( B1 => n11571, B2 => n11557, A => n20354, ZN => 
                           n2781);
   U1514 : AND3_X1 port map( A1 => N114, A2 => n11616, A3 => n11617, ZN => 
                           n11588);
   U1515 : AND3_X1 port map( A1 => N79, A2 => n11565, A3 => n11658, ZN => 
                           n11634);
   U1516 : OAI221_X1 port map( B1 => n1697, B2 => n1726, C1 => n1699, C2 => 
                           n1727, A => n20352, ZN => n1725);
   U1517 : OAI221_X1 port map( B1 => n1697, B2 => n1698, C1 => n1699, C2 => 
                           n1700, A => n20352, ZN => n1633);
   U1518 : OAI221_X1 port map( B1 => n1697, B2 => n1715, C1 => n1699, C2 => 
                           n1716, A => n20352, ZN => n1714);
   U1519 : OAI221_X1 port map( B1 => n1708, B2 => n1726, C1 => n1709, C2 => 
                           n1727, A => n20352, ZN => n1799);
   U1520 : OAI221_X1 port map( B1 => n1708, B2 => n1715, C1 => n1709, C2 => 
                           n1716, A => n20352, ZN => n1721);
   U1521 : OAI221_X1 port map( B1 => n1698, B2 => n1708, C1 => n1700, C2 => 
                           n1709, A => n20352, ZN => n1707);
   U1522 : AND3_X1 port map( A1 => N115, A2 => n11621, A3 => n11617, ZN => 
                           n11590);
   U1523 : AND3_X1 port map( A1 => N80, A2 => n11660, A3 => n11658, ZN => 
                           n11636);
   U1524 : AND3_X1 port map( A1 => N115, A2 => N114, A3 => n11617, ZN => n11594
                           );
   U1525 : AND3_X1 port map( A1 => N80, A2 => N79, A3 => n11658, ZN => n11639);
   U1526 : OAI22_X1 port map( A1 => n2192, A2 => n19171, B1 => n19170, B2 => 
                           n11555, ZN => n11651);
   U1527 : OAI22_X1 port map( A1 => n2192, A2 => n19370, B1 => n19369, B2 => 
                           n11555, ZN => n11610);
   U1528 : OAI22_X1 port map( A1 => n2189, A2 => n19171, B1 => n19170, B2 => 
                           n11487, ZN => n11531);
   U1529 : OAI22_X1 port map( A1 => n2189, A2 => n19370, B1 => n19369, B2 => 
                           n11487, ZN => n11511);
   U1530 : OAI22_X1 port map( A1 => n2186, A2 => n19171, B1 => n19170, B2 => 
                           n11420, ZN => n11464);
   U1531 : OAI22_X1 port map( A1 => n2186, A2 => n19370, B1 => n19369, B2 => 
                           n11420, ZN => n11444);
   U1532 : OAI22_X1 port map( A1 => n2183, A2 => n19171, B1 => n19170, B2 => 
                           n11353, ZN => n11397);
   U1533 : OAI22_X1 port map( A1 => n2183, A2 => n19370, B1 => n19369, B2 => 
                           n11353, ZN => n11376);
   U1534 : OAI22_X1 port map( A1 => n2180, A2 => n19171, B1 => n19170, B2 => 
                           n11286, ZN => n11329);
   U1535 : OAI22_X1 port map( A1 => n2180, A2 => n19370, B1 => n19369, B2 => 
                           n11286, ZN => n11309);
   U1536 : OAI22_X1 port map( A1 => n2177, A2 => n19171, B1 => n19170, B2 => 
                           n11218, ZN => n11262);
   U1537 : OAI22_X1 port map( A1 => n2177, A2 => n19370, B1 => n19369, B2 => 
                           n11218, ZN => n11242);
   U1538 : OAI22_X1 port map( A1 => n2174, A2 => n19171, B1 => n19170, B2 => 
                           n11151, ZN => n11195);
   U1539 : OAI22_X1 port map( A1 => n2174, A2 => n19370, B1 => n19369, B2 => 
                           n11151, ZN => n11175);
   U1540 : OAI22_X1 port map( A1 => n2171, A2 => n19171, B1 => n19170, B2 => 
                           n11084, ZN => n11128);
   U1541 : OAI22_X1 port map( A1 => n2171, A2 => n19370, B1 => n19369, B2 => 
                           n11084, ZN => n11107);
   U1542 : OAI22_X1 port map( A1 => n2168, A2 => n19171, B1 => n19170, B2 => 
                           n11017, ZN => n11060);
   U1543 : OAI22_X1 port map( A1 => n2168, A2 => n19370, B1 => n19369, B2 => 
                           n11017, ZN => n11040);
   U1544 : OAI22_X1 port map( A1 => n2165, A2 => n19171, B1 => n19170, B2 => 
                           n10949, ZN => n10993);
   U1545 : OAI22_X1 port map( A1 => n2165, A2 => n19370, B1 => n19369, B2 => 
                           n10949, ZN => n10973);
   U1546 : OAI22_X1 port map( A1 => n2162, A2 => n19171, B1 => n19170, B2 => 
                           n10882, ZN => n10926);
   U1547 : OAI22_X1 port map( A1 => n2162, A2 => n19370, B1 => n19369, B2 => 
                           n10882, ZN => n10905);
   U1548 : OAI22_X1 port map( A1 => n2159, A2 => n19171, B1 => n19170, B2 => 
                           n10815, ZN => n10859);
   U1549 : OAI22_X1 port map( A1 => n2159, A2 => n19370, B1 => n19369, B2 => 
                           n10815, ZN => n10838);
   U1550 : OAI22_X1 port map( A1 => n2156, A2 => n19172, B1 => n19170, B2 => 
                           n10747, ZN => n10791);
   U1551 : OAI22_X1 port map( A1 => n2156, A2 => n19371, B1 => n19369, B2 => 
                           n10747, ZN => n10771);
   U1552 : OAI22_X1 port map( A1 => n2153, A2 => n19172, B1 => n19169, B2 => 
                           n10680, ZN => n10724);
   U1553 : OAI22_X1 port map( A1 => n2153, A2 => n19371, B1 => n19368, B2 => 
                           n10680, ZN => n10704);
   U1554 : OAI22_X1 port map( A1 => n2150, A2 => n19172, B1 => n19169, B2 => 
                           n10613, ZN => n10657);
   U1555 : OAI22_X1 port map( A1 => n2150, A2 => n19371, B1 => n19368, B2 => 
                           n10613, ZN => n10636);
   U1556 : OAI22_X1 port map( A1 => n2147, A2 => n19172, B1 => n19169, B2 => 
                           n10546, ZN => n10590);
   U1557 : OAI22_X1 port map( A1 => n2147, A2 => n19371, B1 => n19368, B2 => 
                           n10546, ZN => n10569);
   U1558 : OAI22_X1 port map( A1 => n2144, A2 => n19172, B1 => n19169, B2 => 
                           n10478, ZN => n10522);
   U1559 : OAI22_X1 port map( A1 => n2144, A2 => n19371, B1 => n19368, B2 => 
                           n10478, ZN => n10502);
   U1560 : OAI22_X1 port map( A1 => n2143, A2 => n19172, B1 => n19169, B2 => 
                           n10411, ZN => n10455);
   U1561 : OAI22_X1 port map( A1 => n2143, A2 => n19371, B1 => n19368, B2 => 
                           n10411, ZN => n10435);
   U1562 : OAI22_X1 port map( A1 => n2142, A2 => n19172, B1 => n19169, B2 => 
                           n10344, ZN => n10388);
   U1563 : OAI22_X1 port map( A1 => n2142, A2 => n19371, B1 => n19368, B2 => 
                           n10344, ZN => n10367);
   U1564 : OAI22_X1 port map( A1 => n2141, A2 => n19172, B1 => n19169, B2 => 
                           n10277, ZN => n10320);
   U1565 : OAI22_X1 port map( A1 => n2141, A2 => n19371, B1 => n19368, B2 => 
                           n10277, ZN => n10300);
   U1566 : OAI22_X1 port map( A1 => n2140, A2 => n19172, B1 => n19169, B2 => 
                           n10209, ZN => n10253);
   U1567 : OAI22_X1 port map( A1 => n2140, A2 => n19371, B1 => n19368, B2 => 
                           n10209, ZN => n10233);
   U1568 : OAI22_X1 port map( A1 => n2139, A2 => n19172, B1 => n19169, B2 => 
                           n10142, ZN => n10186);
   U1569 : OAI22_X1 port map( A1 => n2139, A2 => n19371, B1 => n19368, B2 => 
                           n10142, ZN => n10166);
   U1570 : OAI22_X1 port map( A1 => n2138, A2 => n19172, B1 => n19169, B2 => 
                           n10075, ZN => n10119);
   U1571 : OAI22_X1 port map( A1 => n2138, A2 => n19371, B1 => n19368, B2 => 
                           n10075, ZN => n10098);
   U1572 : OAI22_X1 port map( A1 => n2137, A2 => n19172, B1 => n19169, B2 => 
                           n10008, ZN => n10051);
   U1573 : OAI22_X1 port map( A1 => n2137, A2 => n19371, B1 => n19368, B2 => 
                           n10008, ZN => n10031);
   U1574 : OAI22_X1 port map( A1 => n2136, A2 => n19173, B1 => n19169, B2 => 
                           n9940, ZN => n9984);
   U1575 : OAI22_X1 port map( A1 => n2136, A2 => n19372, B1 => n19368, B2 => 
                           n9940, ZN => n9964);
   U1576 : OAI22_X1 port map( A1 => n2135, A2 => n19173, B1 => n19169, B2 => 
                           n9873, ZN => n9917);
   U1577 : OAI22_X1 port map( A1 => n2135, A2 => n19372, B1 => n19368, B2 => 
                           n9873, ZN => n9896);
   U1578 : OAI22_X1 port map( A1 => n2134, A2 => n19173, B1 => n19168, B2 => 
                           n9806, ZN => n9850);
   U1579 : OAI22_X1 port map( A1 => n2134, A2 => n19372, B1 => n19367, B2 => 
                           n9806, ZN => n9829);
   U1580 : OAI22_X1 port map( A1 => n2133, A2 => n19173, B1 => n19168, B2 => 
                           n9738, ZN => n9782);
   U1581 : OAI22_X1 port map( A1 => n2133, A2 => n19372, B1 => n19367, B2 => 
                           n9738, ZN => n9762);
   U1582 : OAI22_X1 port map( A1 => n2132, A2 => n19173, B1 => n19168, B2 => 
                           n9671, ZN => n9715);
   U1583 : OAI22_X1 port map( A1 => n2132, A2 => n19372, B1 => n19367, B2 => 
                           n9671, ZN => n9695);
   U1584 : OAI22_X1 port map( A1 => n2131, A2 => n19173, B1 => n19168, B2 => 
                           n9604, ZN => n9648);
   U1585 : OAI22_X1 port map( A1 => n2131, A2 => n19372, B1 => n19367, B2 => 
                           n9604, ZN => n9627);
   U1586 : OAI22_X1 port map( A1 => n2130, A2 => n19173, B1 => n19168, B2 => 
                           n9537, ZN => n9580);
   U1587 : OAI22_X1 port map( A1 => n2130, A2 => n19372, B1 => n19367, B2 => 
                           n9537, ZN => n9560);
   U1588 : OAI22_X1 port map( A1 => n2129, A2 => n19173, B1 => n19168, B2 => 
                           n9469, ZN => n9513);
   U1589 : OAI22_X1 port map( A1 => n2129, A2 => n19372, B1 => n19367, B2 => 
                           n9469, ZN => n9493);
   U1590 : OAI22_X1 port map( A1 => n2128, A2 => n19173, B1 => n19168, B2 => 
                           n9402, ZN => n9446);
   U1591 : OAI22_X1 port map( A1 => n2128, A2 => n19372, B1 => n19367, B2 => 
                           n9402, ZN => n9426);
   U1592 : OAI22_X1 port map( A1 => n2127, A2 => n19173, B1 => n19168, B2 => 
                           n9335, ZN => n9379);
   U1593 : OAI22_X1 port map( A1 => n2127, A2 => n19372, B1 => n19367, B2 => 
                           n9335, ZN => n9358);
   U1594 : OAI22_X1 port map( A1 => n2126, A2 => n19173, B1 => n19168, B2 => 
                           n9268, ZN => n9311);
   U1595 : OAI22_X1 port map( A1 => n2126, A2 => n19372, B1 => n19367, B2 => 
                           n9268, ZN => n9291);
   U1596 : OAI22_X1 port map( A1 => n2125, A2 => n19173, B1 => n19168, B2 => 
                           n6961, ZN => n7004);
   U1597 : OAI22_X1 port map( A1 => n2125, A2 => n19372, B1 => n19367, B2 => 
                           n6961, ZN => n6984);
   U1598 : OAI22_X1 port map( A1 => n2124, A2 => n19174, B1 => n19168, B2 => 
                           n6894, ZN => n6937);
   U1599 : OAI22_X1 port map( A1 => n2124, A2 => n19373, B1 => n19367, B2 => 
                           n6894, ZN => n6917);
   U1600 : OAI22_X1 port map( A1 => n2123, A2 => n19174, B1 => n19168, B2 => 
                           n6827, ZN => n6871);
   U1601 : OAI22_X1 port map( A1 => n2123, A2 => n19373, B1 => n19367, B2 => 
                           n6827, ZN => n6850);
   U1602 : OAI22_X1 port map( A1 => n2122, A2 => n19174, B1 => n19168, B2 => 
                           n6760, ZN => n6804);
   U1603 : OAI22_X1 port map( A1 => n2122, A2 => n19373, B1 => n19367, B2 => 
                           n6760, ZN => n6783);
   U1604 : OAI22_X1 port map( A1 => n2121, A2 => n19174, B1 => n19167, B2 => 
                           n6692, ZN => n6736);
   U1605 : OAI22_X1 port map( A1 => n2121, A2 => n19373, B1 => n19366, B2 => 
                           n6692, ZN => n6716);
   U1606 : OAI22_X1 port map( A1 => n2120, A2 => n19174, B1 => n19167, B2 => 
                           n6625, ZN => n6669);
   U1607 : OAI22_X1 port map( A1 => n2120, A2 => n19373, B1 => n19366, B2 => 
                           n6625, ZN => n6649);
   U1608 : OAI22_X1 port map( A1 => n2119, A2 => n19174, B1 => n19167, B2 => 
                           n6559, ZN => n6602);
   U1609 : OAI22_X1 port map( A1 => n2119, A2 => n19373, B1 => n19366, B2 => 
                           n6559, ZN => n6582);
   U1610 : OAI22_X1 port map( A1 => n2118, A2 => n19174, B1 => n19167, B2 => 
                           n6493, ZN => n6536);
   U1611 : OAI22_X1 port map( A1 => n2118, A2 => n19373, B1 => n19366, B2 => 
                           n6493, ZN => n6516);
   U1612 : OAI22_X1 port map( A1 => n2117, A2 => n19174, B1 => n19167, B2 => 
                           n6427, ZN => n6470);
   U1613 : OAI22_X1 port map( A1 => n2117, A2 => n19373, B1 => n19366, B2 => 
                           n6427, ZN => n6450);
   U1614 : OAI22_X1 port map( A1 => n2116, A2 => n19174, B1 => n19167, B2 => 
                           n6361, ZN => n6404);
   U1615 : OAI22_X1 port map( A1 => n2116, A2 => n19373, B1 => n19366, B2 => 
                           n6361, ZN => n6384);
   U1616 : OAI22_X1 port map( A1 => n2115, A2 => n19174, B1 => n19167, B2 => 
                           n6295, ZN => n6338);
   U1617 : OAI22_X1 port map( A1 => n2115, A2 => n19373, B1 => n19366, B2 => 
                           n6295, ZN => n6318);
   U1618 : OAI22_X1 port map( A1 => n2114, A2 => n19174, B1 => n19167, B2 => 
                           n6229, ZN => n6272);
   U1619 : OAI22_X1 port map( A1 => n2114, A2 => n19373, B1 => n19366, B2 => 
                           n6229, ZN => n6252);
   U1620 : OAI22_X1 port map( A1 => n2113, A2 => n19174, B1 => n19167, B2 => 
                           n6163, ZN => n6206);
   U1621 : OAI22_X1 port map( A1 => n2113, A2 => n19373, B1 => n19366, B2 => 
                           n6163, ZN => n6186);
   U1622 : OAI22_X1 port map( A1 => n2112, A2 => n19175, B1 => n19167, B2 => 
                           n6097, ZN => n6140);
   U1623 : OAI22_X1 port map( A1 => n2112, A2 => n19374, B1 => n19366, B2 => 
                           n6097, ZN => n6120);
   U1624 : OAI22_X1 port map( A1 => n2111, A2 => n19175, B1 => n19167, B2 => 
                           n6029, ZN => n6074);
   U1625 : OAI22_X1 port map( A1 => n2111, A2 => n19374, B1 => n19366, B2 => 
                           n6029, ZN => n6054);
   U1626 : OAI22_X1 port map( A1 => n2110, A2 => n19175, B1 => n19167, B2 => 
                           n5961, ZN => n6006);
   U1627 : OAI22_X1 port map( A1 => n2110, A2 => n19374, B1 => n19366, B2 => 
                           n5961, ZN => n5986);
   U1628 : OAI22_X1 port map( A1 => n2109, A2 => n19175, B1 => n19167, B2 => 
                           n5894, ZN => n5938);
   U1629 : OAI22_X1 port map( A1 => n2109, A2 => n19374, B1 => n19366, B2 => 
                           n5894, ZN => n5918);
   U1630 : OAI22_X1 port map( A1 => n2108, A2 => n19175, B1 => n19166, B2 => 
                           n5827, ZN => n5871);
   U1631 : OAI22_X1 port map( A1 => n2108, A2 => n19374, B1 => n19365, B2 => 
                           n5827, ZN => n5851);
   U1632 : OAI22_X1 port map( A1 => n2107, A2 => n19175, B1 => n19166, B2 => 
                           n5755, ZN => n5804);
   U1633 : OAI22_X1 port map( A1 => n2107, A2 => n19374, B1 => n19365, B2 => 
                           n5755, ZN => n5784);
   U1634 : OAI22_X1 port map( A1 => n2106, A2 => n19175, B1 => n19166, B2 => 
                           n5685, ZN => n5732);
   U1635 : OAI22_X1 port map( A1 => n2106, A2 => n19374, B1 => n19365, B2 => 
                           n5685, ZN => n5712);
   U1636 : OAI22_X1 port map( A1 => n2105, A2 => n19175, B1 => n19166, B2 => 
                           n5617, ZN => n5662);
   U1637 : OAI22_X1 port map( A1 => n2105, A2 => n19374, B1 => n19365, B2 => 
                           n5617, ZN => n5642);
   U1638 : OAI22_X1 port map( A1 => n2104, A2 => n19175, B1 => n19166, B2 => 
                           n5548, ZN => n5594);
   U1639 : OAI22_X1 port map( A1 => n2104, A2 => n19374, B1 => n19365, B2 => 
                           n5548, ZN => n5574);
   U1640 : OAI22_X1 port map( A1 => n2103, A2 => n19175, B1 => n19166, B2 => 
                           n5479, ZN => n5525);
   U1641 : OAI22_X1 port map( A1 => n2103, A2 => n19374, B1 => n19365, B2 => 
                           n5479, ZN => n5505);
   U1642 : OAI22_X1 port map( A1 => n2102, A2 => n19175, B1 => n19166, B2 => 
                           n5411, ZN => n5456);
   U1643 : OAI22_X1 port map( A1 => n2102, A2 => n19374, B1 => n19365, B2 => 
                           n5411, ZN => n5436);
   U1644 : OAI22_X1 port map( A1 => n2101, A2 => n19175, B1 => n19166, B2 => 
                           n5341, ZN => n5388);
   U1645 : OAI22_X1 port map( A1 => n2101, A2 => n19374, B1 => n19365, B2 => 
                           n5341, ZN => n5368);
   U1646 : OAI22_X1 port map( A1 => n2100, A2 => n19176, B1 => n19166, B2 => 
                           n4856, ZN => n5318);
   U1647 : OAI22_X1 port map( A1 => n2100, A2 => n19375, B1 => n19365, B2 => 
                           n4856, ZN => n5298);
   U1648 : OAI22_X1 port map( A1 => n2099, A2 => n19176, B1 => n19166, B2 => 
                           n3638, ZN => n4513);
   U1649 : OAI22_X1 port map( A1 => n2099, A2 => n19375, B1 => n19365, B2 => 
                           n3638, ZN => n4109);
   U1650 : OAI22_X1 port map( A1 => n2098, A2 => n19176, B1 => n19166, B2 => 
                           n3208, ZN => n3294);
   U1651 : OAI22_X1 port map( A1 => n2098, A2 => n19375, B1 => n19365, B2 => 
                           n3208, ZN => n3254);
   U1652 : OAI22_X1 port map( A1 => n2097, A2 => n19176, B1 => n2768, B2 => 
                           n19166, ZN => n3119);
   U1653 : OAI22_X1 port map( A1 => n2097, A2 => n19375, B1 => n2768, B2 => 
                           n19365, ZN => n3002);
   U1654 : NOR3_X1 port map( A1 => n11570, A2 => n11571, A3 => n11572, ZN => 
                           n11569);
   U1655 : XNOR2_X1 port map( A => n1947, B => N114, ZN => n11570);
   U1656 : XNOR2_X1 port map( A => n11573, B => n2228, ZN => n11572);
   U1657 : NAND2_X1 port map( A1 => N149, A2 => n2764, ZN => n2014);
   U1658 : NAND2_X1 port map( A1 => n11684, A2 => n11691, ZN => n3196);
   U1659 : NOR2_X1 port map( A1 => n18915, A2 => n2093, ZN => n11675);
   U1660 : OAI22_X1 port map( A1 => N150, A2 => n11565, B1 => N149, B2 => 
                           n11660, ZN => n11750);
   U1661 : OAI21_X1 port map( B1 => U3_U6_Z_0, B2 => n11748, A => 
                           sub_123_carry_4_port, ZN => n11556);
   U1662 : AOI21_X1 port map( B1 => n11687, B2 => n11681, A => n2086, ZN => 
                           n11715);
   U1663 : INV_X1 port map( A => N148, ZN => n2094);
   U1664 : OAI22_X1 port map( A1 => n2090, A2 => n11694, B1 => n11695, B2 => 
                           n11696, ZN => n11693);
   U1665 : AOI22_X1 port map( A1 => n19183, A2 => n11605, B1 => n19177, B2 => 
                           n11606, ZN => n11646);
   U1666 : AOI22_X1 port map( A1 => n19255, A2 => n11585, B1 => n19249, B2 => 
                           n11586, ZN => n11632);
   U1667 : AOI22_X1 port map( A1 => n19406, A2 => n11598, B1 => n19400, B2 => 
                           n11599, ZN => n11597);
   U1668 : AOI22_X1 port map( A1 => n19454, A2 => n11585, B1 => n19448, B2 => 
                           n11586, ZN => n11584);
   U1669 : AOI22_X1 port map( A1 => n19382, A2 => n11605, B1 => n19376, B2 => 
                           n11606, ZN => n11604);
   U1670 : AOI22_X1 port map( A1 => n19183, A2 => n11506, B1 => n19177, B2 => 
                           n11507, ZN => n11527);
   U1671 : AOI22_X1 port map( A1 => n19255, A2 => n11498, B1 => n19249, B2 => 
                           n11499, ZN => n11524);
   U1672 : AOI22_X1 port map( A1 => n19406, A2 => n11503, B1 => n19400, B2 => 
                           n11504, ZN => n11502);
   U1673 : AOI22_X1 port map( A1 => n19454, A2 => n11498, B1 => n19448, B2 => 
                           n11499, ZN => n11497);
   U1674 : AOI22_X1 port map( A1 => n19382, A2 => n11506, B1 => n19376, B2 => 
                           n11507, ZN => n11505);
   U1675 : AOI22_X1 port map( A1 => n19183, A2 => n11439, B1 => n19177, B2 => 
                           n11440, ZN => n11460);
   U1676 : AOI22_X1 port map( A1 => n19255, A2 => n11430, B1 => n19249, B2 => 
                           n11431, ZN => n11457);
   U1677 : AOI22_X1 port map( A1 => n19406, A2 => n11435, B1 => n19400, B2 => 
                           n11437, ZN => n11434);
   U1678 : AOI22_X1 port map( A1 => n19454, A2 => n11430, B1 => n19448, B2 => 
                           n11431, ZN => n11429);
   U1679 : AOI22_X1 port map( A1 => n19382, A2 => n11439, B1 => n19376, B2 => 
                           n11440, ZN => n11438);
   U1680 : AOI22_X1 port map( A1 => n19183, A2 => n11371, B1 => n19177, B2 => 
                           n11372, ZN => n11393);
   U1681 : AOI22_X1 port map( A1 => n19255, A2 => n11363, B1 => n19249, B2 => 
                           n11364, ZN => n11390);
   U1682 : AOI22_X1 port map( A1 => n19406, A2 => n11368, B1 => n19400, B2 => 
                           n11369, ZN => n11367);
   U1683 : AOI22_X1 port map( A1 => n19454, A2 => n11363, B1 => n19448, B2 => 
                           n11364, ZN => n11362);
   U1684 : AOI22_X1 port map( A1 => n19382, A2 => n11371, B1 => n19376, B2 => 
                           n11372, ZN => n11370);
   U1685 : AOI22_X1 port map( A1 => n19183, A2 => n17722, B1 => n19177, B2 => 
                           n17927, ZN => n11325);
   U1686 : AOI22_X1 port map( A1 => n19255, A2 => n17936, B1 => n19249, B2 => 
                           n17807, ZN => n11322);
   U1687 : AOI22_X1 port map( A1 => n19406, A2 => n17868, B1 => n19400, B2 => 
                           n18108, ZN => n11300);
   U1688 : AOI22_X1 port map( A1 => n19454, A2 => n17936, B1 => n19448, B2 => 
                           n17807, ZN => n11295);
   U1689 : AOI22_X1 port map( A1 => n19382, A2 => n17722, B1 => n19376, B2 => 
                           n17927, ZN => n11303);
   U1690 : AOI22_X1 port map( A1 => n19183, A2 => n17723, B1 => n19177, B2 => 
                           n17928, ZN => n11258);
   U1691 : AOI22_X1 port map( A1 => n19255, A2 => n17937, B1 => n19249, B2 => 
                           n17808, ZN => n11255);
   U1692 : AOI22_X1 port map( A1 => n19406, A2 => n17869, B1 => n19400, B2 => 
                           n18109, ZN => n11233);
   U1693 : AOI22_X1 port map( A1 => n19454, A2 => n17937, B1 => n19448, B2 => 
                           n17808, ZN => n11228);
   U1694 : AOI22_X1 port map( A1 => n19382, A2 => n17723, B1 => n19376, B2 => 
                           n17928, ZN => n11236);
   U1695 : AOI22_X1 port map( A1 => n19183, A2 => n17724, B1 => n19177, B2 => 
                           n17929, ZN => n11191);
   U1696 : AOI22_X1 port map( A1 => n19255, A2 => n17938, B1 => n19249, B2 => 
                           n17809, ZN => n11188);
   U1697 : AOI22_X1 port map( A1 => n19406, A2 => n17870, B1 => n19400, B2 => 
                           n18110, ZN => n11165);
   U1698 : AOI22_X1 port map( A1 => n19454, A2 => n17938, B1 => n19448, B2 => 
                           n17809, ZN => n11160);
   U1699 : AOI22_X1 port map( A1 => n19382, A2 => n17724, B1 => n19376, B2 => 
                           n17929, ZN => n11168);
   U1700 : AOI22_X1 port map( A1 => n19183, A2 => n17725, B1 => n19177, B2 => 
                           n17930, ZN => n11124);
   U1701 : AOI22_X1 port map( A1 => n19255, A2 => n17939, B1 => n19249, B2 => 
                           n17810, ZN => n11121);
   U1702 : AOI22_X1 port map( A1 => n19406, A2 => n17871, B1 => n19400, B2 => 
                           n18111, ZN => n11098);
   U1703 : AOI22_X1 port map( A1 => n19454, A2 => n17939, B1 => n19448, B2 => 
                           n17810, ZN => n11093);
   U1704 : AOI22_X1 port map( A1 => n19382, A2 => n17725, B1 => n19376, B2 => 
                           n17930, ZN => n11101);
   U1705 : AOI22_X1 port map( A1 => n19183, A2 => n17726, B1 => n19177, B2 => 
                           n17931, ZN => n11056);
   U1706 : AOI22_X1 port map( A1 => n19255, A2 => n17940, B1 => n19249, B2 => 
                           n17811, ZN => n11053);
   U1707 : AOI22_X1 port map( A1 => n19406, A2 => n17872, B1 => n19400, B2 => 
                           n18112, ZN => n11031);
   U1708 : AOI22_X1 port map( A1 => n19454, A2 => n17940, B1 => n19448, B2 => 
                           n17811, ZN => n11026);
   U1709 : AOI22_X1 port map( A1 => n19382, A2 => n17726, B1 => n19376, B2 => 
                           n17931, ZN => n11034);
   U1710 : AOI22_X1 port map( A1 => n19183, A2 => n17727, B1 => n19177, B2 => 
                           n17932, ZN => n10989);
   U1711 : AOI22_X1 port map( A1 => n19255, A2 => n17941, B1 => n19249, B2 => 
                           n17812, ZN => n10986);
   U1712 : AOI22_X1 port map( A1 => n19406, A2 => n17873, B1 => n19400, B2 => 
                           n18113, ZN => n10964);
   U1713 : AOI22_X1 port map( A1 => n19454, A2 => n17941, B1 => n19448, B2 => 
                           n17812, ZN => n10958);
   U1714 : AOI22_X1 port map( A1 => n19382, A2 => n17727, B1 => n19376, B2 => 
                           n17932, ZN => n10967);
   U1715 : AOI22_X1 port map( A1 => n19183, A2 => n17728, B1 => n19177, B2 => 
                           n17933, ZN => n10922);
   U1716 : AOI22_X1 port map( A1 => n19255, A2 => n17942, B1 => n19249, B2 => 
                           n17813, ZN => n10919);
   U1717 : AOI22_X1 port map( A1 => n19406, A2 => n17874, B1 => n19400, B2 => 
                           n18114, ZN => n10896);
   U1718 : AOI22_X1 port map( A1 => n19454, A2 => n17942, B1 => n19448, B2 => 
                           n17813, ZN => n10891);
   U1719 : AOI22_X1 port map( A1 => n19382, A2 => n17728, B1 => n19376, B2 => 
                           n17933, ZN => n10899);
   U1720 : AOI22_X1 port map( A1 => n19183, A2 => n17729, B1 => n19177, B2 => 
                           n17934, ZN => n10855);
   U1721 : AOI22_X1 port map( A1 => n19255, A2 => n17943, B1 => n19249, B2 => 
                           n17814, ZN => n10851);
   U1722 : AOI22_X1 port map( A1 => n19406, A2 => n17875, B1 => n19400, B2 => 
                           n18115, ZN => n10829);
   U1723 : AOI22_X1 port map( A1 => n19454, A2 => n17943, B1 => n19448, B2 => 
                           n17814, ZN => n10824);
   U1724 : AOI22_X1 port map( A1 => n19382, A2 => n17729, B1 => n19376, B2 => 
                           n17934, ZN => n10832);
   U1726 : AOI22_X1 port map( A1 => n19184, A2 => n17730, B1 => n19178, B2 => 
                           n17888, ZN => n10787);
   U1727 : AOI22_X1 port map( A1 => n19256, A2 => n17944, B1 => n19250, B2 => 
                           n17768, ZN => n10784);
   U1728 : AOI22_X1 port map( A1 => n19407, A2 => n17816, B1 => n19401, B2 => 
                           n18056, ZN => n10762);
   U1729 : AOI22_X1 port map( A1 => n19455, A2 => n17944, B1 => n19449, B2 => 
                           n17768, ZN => n10757);
   U1730 : AOI22_X1 port map( A1 => n19383, A2 => n17730, B1 => n19377, B2 => 
                           n17888, ZN => n10765);
   U1731 : AOI22_X1 port map( A1 => n19184, A2 => n17731, B1 => n19178, B2 => 
                           n17889, ZN => n10720);
   U1732 : AOI22_X1 port map( A1 => n19256, A2 => n17945, B1 => n19250, B2 => 
                           n17769, ZN => n10717);
   U1733 : AOI22_X1 port map( A1 => n19407, A2 => n17817, B1 => n19401, B2 => 
                           n18057, ZN => n10694);
   U1734 : AOI22_X1 port map( A1 => n19455, A2 => n17945, B1 => n19449, B2 => 
                           n17769, ZN => n10689);
   U1735 : AOI22_X1 port map( A1 => n19383, A2 => n17731, B1 => n19377, B2 => 
                           n17889, ZN => n10698);
   U1736 : AOI22_X1 port map( A1 => n19184, A2 => n17732, B1 => n19178, B2 => 
                           n17890, ZN => n10653);
   U1737 : AOI22_X1 port map( A1 => n19256, A2 => n17946, B1 => n19250, B2 => 
                           n17770, ZN => n10650);
   U1738 : AOI22_X1 port map( A1 => n19407, A2 => n17818, B1 => n19401, B2 => 
                           n18058, ZN => n10627);
   U1739 : AOI22_X1 port map( A1 => n19455, A2 => n17946, B1 => n19449, B2 => 
                           n17770, ZN => n10622);
   U1740 : AOI22_X1 port map( A1 => n19383, A2 => n17732, B1 => n19377, B2 => 
                           n17890, ZN => n10630);
   U1741 : AOI22_X1 port map( A1 => n19184, A2 => n17733, B1 => n19178, B2 => 
                           n17891, ZN => n10585);
   U1742 : AOI22_X1 port map( A1 => n19256, A2 => n17947, B1 => n19250, B2 => 
                           n17771, ZN => n10582);
   U1743 : AOI22_X1 port map( A1 => n19407, A2 => n17819, B1 => n19401, B2 => 
                           n18059, ZN => n10560);
   U1744 : AOI22_X1 port map( A1 => n19455, A2 => n17947, B1 => n19449, B2 => 
                           n17771, ZN => n10555);
   U1745 : AOI22_X1 port map( A1 => n19383, A2 => n17733, B1 => n19377, B2 => 
                           n17891, ZN => n10563);
   U1746 : AOI22_X1 port map( A1 => n19184, A2 => n17734, B1 => n19178, B2 => 
                           n17892, ZN => n10518);
   U1747 : AOI22_X1 port map( A1 => n19256, A2 => n17948, B1 => n19250, B2 => 
                           n17772, ZN => n10515);
   U1748 : AOI22_X1 port map( A1 => n19407, A2 => n17820, B1 => n19401, B2 => 
                           n18060, ZN => n10493);
   U1749 : AOI22_X1 port map( A1 => n19455, A2 => n17948, B1 => n19449, B2 => 
                           n17772, ZN => n10488);
   U1750 : AOI22_X1 port map( A1 => n19383, A2 => n17734, B1 => n19377, B2 => 
                           n17892, ZN => n10496);
   U1751 : AOI22_X1 port map( A1 => n19184, A2 => n17735, B1 => n19178, B2 => 
                           n17893, ZN => n10451);
   U1752 : AOI22_X1 port map( A1 => n19256, A2 => n17949, B1 => n19250, B2 => 
                           n17773, ZN => n10448);
   U1753 : AOI22_X1 port map( A1 => n19407, A2 => n17821, B1 => n19401, B2 => 
                           n18061, ZN => n10425);
   U1754 : AOI22_X1 port map( A1 => n19455, A2 => n17949, B1 => n19449, B2 => 
                           n17773, ZN => n10420);
   U1755 : AOI22_X1 port map( A1 => n19383, A2 => n17735, B1 => n19377, B2 => 
                           n17893, ZN => n10428);
   U1756 : AOI22_X1 port map( A1 => n19184, A2 => n17736, B1 => n19178, B2 => 
                           n17894, ZN => n10384);
   U1757 : AOI22_X1 port map( A1 => n19256, A2 => n17950, B1 => n19250, B2 => 
                           n17774, ZN => n10381);
   U1758 : AOI22_X1 port map( A1 => n19407, A2 => n17822, B1 => n19401, B2 => 
                           n18062, ZN => n10358);
   U1759 : AOI22_X1 port map( A1 => n19455, A2 => n17950, B1 => n19449, B2 => 
                           n17774, ZN => n10353);
   U1760 : AOI22_X1 port map( A1 => n19383, A2 => n17736, B1 => n19377, B2 => 
                           n17894, ZN => n10361);
   U1761 : AOI22_X1 port map( A1 => n19184, A2 => n17737, B1 => n19178, B2 => 
                           n17895, ZN => n10316);
   U1762 : AOI22_X1 port map( A1 => n19256, A2 => n17951, B1 => n19250, B2 => 
                           n17775, ZN => n10313);
   U1763 : AOI22_X1 port map( A1 => n19407, A2 => n17823, B1 => n19401, B2 => 
                           n18063, ZN => n10291);
   U1764 : AOI22_X1 port map( A1 => n19455, A2 => n17951, B1 => n19449, B2 => 
                           n17775, ZN => n10286);
   U1765 : AOI22_X1 port map( A1 => n19383, A2 => n17737, B1 => n19377, B2 => 
                           n17895, ZN => n10294);
   U1766 : AOI22_X1 port map( A1 => n19184, A2 => n17738, B1 => n19178, B2 => 
                           n17896, ZN => n10249);
   U1767 : AOI22_X1 port map( A1 => n19256, A2 => n17952, B1 => n19250, B2 => 
                           n17776, ZN => n10246);
   U1768 : AOI22_X1 port map( A1 => n19407, A2 => n17824, B1 => n19401, B2 => 
                           n18064, ZN => n10224);
   U1769 : AOI22_X1 port map( A1 => n19455, A2 => n17952, B1 => n19449, B2 => 
                           n17776, ZN => n10219);
   U1770 : AOI22_X1 port map( A1 => n19383, A2 => n17738, B1 => n19377, B2 => 
                           n17896, ZN => n10227);
   U1771 : AOI22_X1 port map( A1 => n19184, A2 => n17739, B1 => n19178, B2 => 
                           n17897, ZN => n10182);
   U1772 : AOI22_X1 port map( A1 => n19256, A2 => n17953, B1 => n19250, B2 => 
                           n17777, ZN => n10179);
   U1773 : AOI22_X1 port map( A1 => n19407, A2 => n17825, B1 => n19401, B2 => 
                           n18065, ZN => n10156);
   U1774 : AOI22_X1 port map( A1 => n19455, A2 => n17953, B1 => n19449, B2 => 
                           n17777, ZN => n10151);
   U1775 : AOI22_X1 port map( A1 => n19383, A2 => n17739, B1 => n19377, B2 => 
                           n17897, ZN => n10159);
   U1776 : AOI22_X1 port map( A1 => n19184, A2 => n17740, B1 => n19178, B2 => 
                           n17898, ZN => n10115);
   U1777 : AOI22_X1 port map( A1 => n19256, A2 => n17954, B1 => n19250, B2 => 
                           n17778, ZN => n10111);
   U1778 : AOI22_X1 port map( A1 => n19407, A2 => n17826, B1 => n19401, B2 => 
                           n18066, ZN => n10089);
   U1779 : AOI22_X1 port map( A1 => n19455, A2 => n17954, B1 => n19449, B2 => 
                           n17778, ZN => n10084);
   U1780 : AOI22_X1 port map( A1 => n19383, A2 => n17740, B1 => n19377, B2 => 
                           n17898, ZN => n10092);
   U1781 : AOI22_X1 port map( A1 => n19184, A2 => n17741, B1 => n19178, B2 => 
                           n17899, ZN => n10047);
   U1782 : AOI22_X1 port map( A1 => n19256, A2 => n17955, B1 => n19250, B2 => 
                           n17779, ZN => n10044);
   U1783 : AOI22_X1 port map( A1 => n19407, A2 => n17827, B1 => n19401, B2 => 
                           n18067, ZN => n10022);
   U1784 : AOI22_X1 port map( A1 => n19455, A2 => n17955, B1 => n19449, B2 => 
                           n17779, ZN => n10017);
   U1785 : AOI22_X1 port map( A1 => n19383, A2 => n17741, B1 => n19377, B2 => 
                           n17899, ZN => n10025);
   U1786 : AOI22_X1 port map( A1 => n19185, A2 => n17742, B1 => n19179, B2 => 
                           n17900, ZN => n9980);
   U1787 : AOI22_X1 port map( A1 => n19257, A2 => n17956, B1 => n19251, B2 => 
                           n17780, ZN => n9977);
   U1788 : AOI22_X1 port map( A1 => n19408, A2 => n17828, B1 => n19402, B2 => 
                           n18068, ZN => n9955);
   U1789 : AOI22_X1 port map( A1 => n19456, A2 => n17956, B1 => n19450, B2 => 
                           n17780, ZN => n9949);
   U1790 : AOI22_X1 port map( A1 => n19384, A2 => n17742, B1 => n19378, B2 => 
                           n17900, ZN => n9958);
   U1791 : AOI22_X1 port map( A1 => n19185, A2 => n17743, B1 => n19179, B2 => 
                           n17901, ZN => n9913);
   U1792 : AOI22_X1 port map( A1 => n19257, A2 => n17957, B1 => n19251, B2 => 
                           n17781, ZN => n9910);
   U1793 : AOI22_X1 port map( A1 => n19408, A2 => n17829, B1 => n19402, B2 => 
                           n18069, ZN => n9887);
   U1794 : AOI22_X1 port map( A1 => n19456, A2 => n17957, B1 => n19450, B2 => 
                           n17781, ZN => n9882);
   U1795 : AOI22_X1 port map( A1 => n19384, A2 => n17743, B1 => n19378, B2 => 
                           n17901, ZN => n9890);
   U1796 : AOI22_X1 port map( A1 => n19185, A2 => n17744, B1 => n19179, B2 => 
                           n17902, ZN => n9845);
   U1797 : AOI22_X1 port map( A1 => n19257, A2 => n17958, B1 => n19251, B2 => 
                           n17782, ZN => n9842);
   U1798 : AOI22_X1 port map( A1 => n19408, A2 => n17830, B1 => n19402, B2 => 
                           n18070, ZN => n9820);
   U1799 : AOI22_X1 port map( A1 => n19456, A2 => n17958, B1 => n19450, B2 => 
                           n17782, ZN => n9815);
   U1800 : AOI22_X1 port map( A1 => n19384, A2 => n17744, B1 => n19378, B2 => 
                           n17902, ZN => n9823);
   U1801 : AOI22_X1 port map( A1 => n19185, A2 => n17745, B1 => n19179, B2 => 
                           n17903, ZN => n9778);
   U1802 : AOI22_X1 port map( A1 => n19257, A2 => n17959, B1 => n19251, B2 => 
                           n17783, ZN => n9775);
   U1803 : AOI22_X1 port map( A1 => n19408, A2 => n17831, B1 => n19402, B2 => 
                           n18071, ZN => n9753);
   U1804 : AOI22_X1 port map( A1 => n19456, A2 => n17959, B1 => n19450, B2 => 
                           n17783, ZN => n9748);
   U1805 : AOI22_X1 port map( A1 => n19384, A2 => n17745, B1 => n19378, B2 => 
                           n17903, ZN => n9756);
   U1806 : AOI22_X1 port map( A1 => n19185, A2 => n17746, B1 => n19179, B2 => 
                           n17904, ZN => n9711);
   U1807 : AOI22_X1 port map( A1 => n19257, A2 => n17960, B1 => n19251, B2 => 
                           n17784, ZN => n9708);
   U1808 : AOI22_X1 port map( A1 => n19408, A2 => n17832, B1 => n19402, B2 => 
                           n18072, ZN => n9685);
   U1809 : AOI22_X1 port map( A1 => n19456, A2 => n17960, B1 => n19450, B2 => 
                           n17784, ZN => n9680);
   U1810 : AOI22_X1 port map( A1 => n19384, A2 => n17746, B1 => n19378, B2 => 
                           n17904, ZN => n9688);
   U1811 : AOI22_X1 port map( A1 => n19185, A2 => n17747, B1 => n19179, B2 => 
                           n17905, ZN => n9644);
   U1812 : AOI22_X1 port map( A1 => n19257, A2 => n17961, B1 => n19251, B2 => 
                           n17785, ZN => n9641);
   U1813 : AOI22_X1 port map( A1 => n19408, A2 => n17833, B1 => n19402, B2 => 
                           n18073, ZN => n9618);
   U1814 : AOI22_X1 port map( A1 => n19456, A2 => n17961, B1 => n19450, B2 => 
                           n17785, ZN => n9613);
   U1815 : AOI22_X1 port map( A1 => n19384, A2 => n17747, B1 => n19378, B2 => 
                           n17905, ZN => n9621);
   U1816 : AOI22_X1 port map( A1 => n19185, A2 => n17748, B1 => n19179, B2 => 
                           n17906, ZN => n9576);
   U1817 : AOI22_X1 port map( A1 => n19257, A2 => n17962, B1 => n19251, B2 => 
                           n17786, ZN => n9573);
   U1818 : AOI22_X1 port map( A1 => n19408, A2 => n17834, B1 => n19402, B2 => 
                           n18074, ZN => n9551);
   U1819 : AOI22_X1 port map( A1 => n19456, A2 => n17962, B1 => n19450, B2 => 
                           n17786, ZN => n9546);
   U1820 : AOI22_X1 port map( A1 => n19384, A2 => n17748, B1 => n19378, B2 => 
                           n17906, ZN => n9554);
   U1821 : AOI22_X1 port map( A1 => n19185, A2 => n17749, B1 => n19179, B2 => 
                           n17907, ZN => n9509);
   U1822 : AOI22_X1 port map( A1 => n19257, A2 => n17963, B1 => n19251, B2 => 
                           n17787, ZN => n9506);
   U1823 : AOI22_X1 port map( A1 => n19408, A2 => n17835, B1 => n19402, B2 => 
                           n18075, ZN => n9484);
   U1824 : AOI22_X1 port map( A1 => n19456, A2 => n17963, B1 => n19450, B2 => 
                           n17787, ZN => n9479);
   U1825 : AOI22_X1 port map( A1 => n19384, A2 => n17749, B1 => n19378, B2 => 
                           n17907, ZN => n9487);
   U1826 : AOI22_X1 port map( A1 => n19185, A2 => n17750, B1 => n19179, B2 => 
                           n17908, ZN => n9442);
   U1827 : AOI22_X1 port map( A1 => n19257, A2 => n17964, B1 => n19251, B2 => 
                           n17788, ZN => n9439);
   U1828 : AOI22_X1 port map( A1 => n19408, A2 => n17836, B1 => n19402, B2 => 
                           n18076, ZN => n9416);
   U1829 : AOI22_X1 port map( A1 => n19456, A2 => n17964, B1 => n19450, B2 => 
                           n17788, ZN => n9411);
   U1830 : AOI22_X1 port map( A1 => n19384, A2 => n17750, B1 => n19378, B2 => 
                           n17908, ZN => n9419);
   U1831 : AOI22_X1 port map( A1 => n19185, A2 => n17751, B1 => n19179, B2 => 
                           n17909, ZN => n9375);
   U1832 : AOI22_X1 port map( A1 => n19257, A2 => n17965, B1 => n19251, B2 => 
                           n17789, ZN => n9372);
   U1833 : AOI22_X1 port map( A1 => n19408, A2 => n17837, B1 => n19402, B2 => 
                           n18077, ZN => n9349);
   U1834 : AOI22_X1 port map( A1 => n19456, A2 => n17965, B1 => n19450, B2 => 
                           n17789, ZN => n9344);
   U1835 : AOI22_X1 port map( A1 => n19384, A2 => n17751, B1 => n19378, B2 => 
                           n17909, ZN => n9352);
   U1836 : AOI22_X1 port map( A1 => n19185, A2 => n17752, B1 => n19179, B2 => 
                           n17910, ZN => n9307);
   U1837 : AOI22_X1 port map( A1 => n19257, A2 => n17966, B1 => n19251, B2 => 
                           n17790, ZN => n9304);
   U1838 : AOI22_X1 port map( A1 => n19408, A2 => n17838, B1 => n19402, B2 => 
                           n18078, ZN => n9282);
   U1839 : AOI22_X1 port map( A1 => n19456, A2 => n17966, B1 => n19450, B2 => 
                           n17790, ZN => n9277);
   U1840 : AOI22_X1 port map( A1 => n19384, A2 => n17752, B1 => n19378, B2 => 
                           n17910, ZN => n9285);
   U1841 : AOI22_X1 port map( A1 => n19185, A2 => n17753, B1 => n19179, B2 => 
                           n17911, ZN => n7000);
   U1842 : AOI22_X1 port map( A1 => n19257, A2 => n17967, B1 => n19251, B2 => 
                           n17791, ZN => n6997);
   U1843 : AOI22_X1 port map( A1 => n19408, A2 => n17839, B1 => n19402, B2 => 
                           n18079, ZN => n6975);
   U1844 : AOI22_X1 port map( A1 => n19456, A2 => n17967, B1 => n19450, B2 => 
                           n17791, ZN => n6970);
   U1845 : AOI22_X1 port map( A1 => n19384, A2 => n17753, B1 => n19378, B2 => 
                           n17911, ZN => n6978);
   U1846 : AOI22_X1 port map( A1 => n19186, A2 => n17754, B1 => n19180, B2 => 
                           n17925, ZN => n6933);
   U1847 : AOI22_X1 port map( A1 => n19258, A2 => n17968, B1 => n19252, B2 => 
                           n17805, ZN => n6930);
   U1848 : AOI22_X1 port map( A1 => n19409, A2 => n17840, B1 => n19403, B2 => 
                           n18080, ZN => n6908);
   U1849 : AOI22_X1 port map( A1 => n19457, A2 => n17968, B1 => n19451, B2 => 
                           n17805, ZN => n6903);
   U1850 : AOI22_X1 port map( A1 => n19385, A2 => n17754, B1 => n19379, B2 => 
                           n17925, ZN => n6911);
   U1851 : AOI22_X1 port map( A1 => n19186, A2 => n17755, B1 => n19180, B2 => 
                           n17926, ZN => n6866);
   U1852 : AOI22_X1 port map( A1 => n19258, A2 => n17969, B1 => n19252, B2 => 
                           n17806, ZN => n6863);
   U1853 : AOI22_X1 port map( A1 => n19409, A2 => n17841, B1 => n19403, B2 => 
                           n18081, ZN => n6841);
   U1854 : AOI22_X1 port map( A1 => n19457, A2 => n17969, B1 => n19451, B2 => 
                           n17806, ZN => n6836);
   U1855 : AOI22_X1 port map( A1 => n19385, A2 => n17755, B1 => n19379, B2 => 
                           n17926, ZN => n6844);
   U1856 : AOI22_X1 port map( A1 => n19186, A2 => n17696, B1 => n19180, B2 => 
                           n17935, ZN => n6799);
   U1857 : AOI22_X1 port map( A1 => n19258, A2 => n17970, B1 => n19252, B2 => 
                           n17815, ZN => n6796);
   U1858 : AOI22_X1 port map( A1 => n19409, A2 => n17842, B1 => n19403, B2 => 
                           n18082, ZN => n6774);
   U1859 : AOI22_X1 port map( A1 => n19457, A2 => n17970, B1 => n19451, B2 => 
                           n17815, ZN => n6769);
   U1860 : AOI22_X1 port map( A1 => n19385, A2 => n17696, B1 => n19379, B2 => 
                           n17935, ZN => n6777);
   U1861 : AOI22_X1 port map( A1 => n19186, A2 => n17701, B1 => n19180, B2 => 
                           n17916, ZN => n6732);
   U1862 : AOI22_X1 port map( A1 => n19258, A2 => n17971, B1 => n19252, B2 => 
                           n17796, ZN => n6729);
   U1863 : AOI22_X1 port map( A1 => n19409, A2 => n17843, B1 => n19403, B2 => 
                           n18083, ZN => n6707);
   U1864 : AOI22_X1 port map( A1 => n19457, A2 => n17971, B1 => n19451, B2 => 
                           n17796, ZN => n6702);
   U1865 : AOI22_X1 port map( A1 => n19385, A2 => n17701, B1 => n19379, B2 => 
                           n17916, ZN => n6710);
   U1866 : AOI22_X1 port map( A1 => n19186, A2 => n17702, B1 => n19180, B2 => 
                           n17917, ZN => n6665);
   U1867 : AOI22_X1 port map( A1 => n19258, A2 => n17972, B1 => n19252, B2 => 
                           n17797, ZN => n6662);
   U1868 : AOI22_X1 port map( A1 => n19409, A2 => n17844, B1 => n19403, B2 => 
                           n18084, ZN => n6639);
   U1869 : AOI22_X1 port map( A1 => n19457, A2 => n17972, B1 => n19451, B2 => 
                           n17797, ZN => n6634);
   U1870 : AOI22_X1 port map( A1 => n19385, A2 => n17702, B1 => n19379, B2 => 
                           n17917, ZN => n6642);
   U1871 : AOI22_X1 port map( A1 => n19186, A2 => n17703, B1 => n19180, B2 => 
                           n17918, ZN => n6598);
   U1872 : AOI22_X1 port map( A1 => n19258, A2 => n17973, B1 => n19252, B2 => 
                           n17798, ZN => n6595);
   U1873 : AOI22_X1 port map( A1 => n19409, A2 => n17845, B1 => n19403, B2 => 
                           n18085, ZN => n6573);
   U1874 : AOI22_X1 port map( A1 => n19457, A2 => n17973, B1 => n19451, B2 => 
                           n17798, ZN => n6568);
   U1875 : AOI22_X1 port map( A1 => n19385, A2 => n17703, B1 => n19379, B2 => 
                           n17918, ZN => n6576);
   U1876 : AOI22_X1 port map( A1 => n19186, A2 => n17704, B1 => n19180, B2 => 
                           n17919, ZN => n6532);
   U1877 : AOI22_X1 port map( A1 => n19258, A2 => n17974, B1 => n19252, B2 => 
                           n17799, ZN => n6529);
   U1878 : AOI22_X1 port map( A1 => n19409, A2 => n17846, B1 => n19403, B2 => 
                           n18086, ZN => n6507);
   U1879 : AOI22_X1 port map( A1 => n19457, A2 => n17974, B1 => n19451, B2 => 
                           n17799, ZN => n6502);
   U1880 : AOI22_X1 port map( A1 => n19385, A2 => n17704, B1 => n19379, B2 => 
                           n17919, ZN => n6510);
   U1881 : AOI22_X1 port map( A1 => n19186, A2 => n17705, B1 => n19180, B2 => 
                           n17920, ZN => n6466);
   U1882 : AOI22_X1 port map( A1 => n19258, A2 => n17975, B1 => n19252, B2 => 
                           n17800, ZN => n6463);
   U1883 : AOI22_X1 port map( A1 => n19409, A2 => n17847, B1 => n19403, B2 => 
                           n18087, ZN => n6441);
   U1884 : AOI22_X1 port map( A1 => n19457, A2 => n17975, B1 => n19451, B2 => 
                           n17800, ZN => n6436);
   U1885 : AOI22_X1 port map( A1 => n19385, A2 => n17705, B1 => n19379, B2 => 
                           n17920, ZN => n6444);
   U1886 : AOI22_X1 port map( A1 => n19186, A2 => n17706, B1 => n19180, B2 => 
                           n17921, ZN => n6400);
   U1887 : AOI22_X1 port map( A1 => n19258, A2 => n17976, B1 => n19252, B2 => 
                           n17801, ZN => n6397);
   U1888 : AOI22_X1 port map( A1 => n19409, A2 => n17848, B1 => n19403, B2 => 
                           n18088, ZN => n6375);
   U1889 : AOI22_X1 port map( A1 => n19457, A2 => n17976, B1 => n19451, B2 => 
                           n17801, ZN => n6370);
   U1890 : AOI22_X1 port map( A1 => n19385, A2 => n17706, B1 => n19379, B2 => 
                           n17921, ZN => n6378);
   U1891 : AOI22_X1 port map( A1 => n19186, A2 => n17707, B1 => n19180, B2 => 
                           n17922, ZN => n6334);
   U1892 : AOI22_X1 port map( A1 => n19258, A2 => n17977, B1 => n19252, B2 => 
                           n17802, ZN => n6331);
   U1893 : AOI22_X1 port map( A1 => n19409, A2 => n17849, B1 => n19403, B2 => 
                           n18089, ZN => n6309);
   U1894 : AOI22_X1 port map( A1 => n19457, A2 => n17977, B1 => n19451, B2 => 
                           n17802, ZN => n6304);
   U1895 : AOI22_X1 port map( A1 => n19385, A2 => n17707, B1 => n19379, B2 => 
                           n17922, ZN => n6312);
   U1896 : AOI22_X1 port map( A1 => n19186, A2 => n17708, B1 => n19180, B2 => 
                           n17923, ZN => n6268);
   U1897 : AOI22_X1 port map( A1 => n19258, A2 => n17978, B1 => n19252, B2 => 
                           n17803, ZN => n6265);
   U1898 : AOI22_X1 port map( A1 => n19409, A2 => n17850, B1 => n19403, B2 => 
                           n18090, ZN => n6243);
   U1899 : AOI22_X1 port map( A1 => n19457, A2 => n17978, B1 => n19451, B2 => 
                           n17803, ZN => n6238);
   U1900 : AOI22_X1 port map( A1 => n19385, A2 => n17708, B1 => n19379, B2 => 
                           n17923, ZN => n6246);
   U1901 : AOI22_X1 port map( A1 => n19186, A2 => n17709, B1 => n19180, B2 => 
                           n17924, ZN => n6202);
   U1902 : AOI22_X1 port map( A1 => n19258, A2 => n17979, B1 => n19252, B2 => 
                           n17804, ZN => n6199);
   U1903 : AOI22_X1 port map( A1 => n19409, A2 => n17851, B1 => n19403, B2 => 
                           n18091, ZN => n6177);
   U1904 : AOI22_X1 port map( A1 => n19457, A2 => n17979, B1 => n19451, B2 => 
                           n17804, ZN => n6172);
   U1905 : AOI22_X1 port map( A1 => n19385, A2 => n17709, B1 => n19379, B2 => 
                           n17924, ZN => n6180);
   U1906 : AOI22_X1 port map( A1 => n19187, A2 => n17710, B1 => n19181, B2 => 
                           n17876, ZN => n6136);
   U1907 : AOI22_X1 port map( A1 => n19259, A2 => n17980, B1 => n19253, B2 => 
                           n17756, ZN => n6133);
   U1908 : AOI22_X1 port map( A1 => n19410, A2 => n17852, B1 => n19404, B2 => 
                           n18092, ZN => n6111);
   U1909 : AOI22_X1 port map( A1 => n19458, A2 => n17980, B1 => n19452, B2 => 
                           n17756, ZN => n6106);
   U1910 : AOI22_X1 port map( A1 => n19386, A2 => n17710, B1 => n19380, B2 => 
                           n17876, ZN => n6114);
   U1911 : AOI22_X1 port map( A1 => n19187, A2 => n17711, B1 => n19181, B2 => 
                           n17877, ZN => n6070);
   U1912 : AOI22_X1 port map( A1 => n19259, A2 => n17981, B1 => n19253, B2 => 
                           n17757, ZN => n6067);
   U1913 : AOI22_X1 port map( A1 => n19410, A2 => n17853, B1 => n19404, B2 => 
                           n18093, ZN => n6045);
   U1914 : AOI22_X1 port map( A1 => n19458, A2 => n17981, B1 => n19452, B2 => 
                           n17757, ZN => n6040);
   U1915 : AOI22_X1 port map( A1 => n19386, A2 => n17711, B1 => n19380, B2 => 
                           n17877, ZN => n6048);
   U1916 : AOI22_X1 port map( A1 => n19187, A2 => n17712, B1 => n19181, B2 => 
                           n17878, ZN => n6002);
   U1917 : AOI22_X1 port map( A1 => n19259, A2 => n17982, B1 => n19253, B2 => 
                           n17758, ZN => n5999);
   U1918 : AOI22_X1 port map( A1 => n19410, A2 => n17854, B1 => n19404, B2 => 
                           n18094, ZN => n5977);
   U1919 : AOI22_X1 port map( A1 => n19458, A2 => n17982, B1 => n19452, B2 => 
                           n17758, ZN => n5972);
   U1920 : AOI22_X1 port map( A1 => n19386, A2 => n17712, B1 => n19380, B2 => 
                           n17878, ZN => n5980);
   U1921 : AOI22_X1 port map( A1 => n19187, A2 => n17713, B1 => n19181, B2 => 
                           n17879, ZN => n5934);
   U1922 : AOI22_X1 port map( A1 => n19259, A2 => n17983, B1 => n19253, B2 => 
                           n17759, ZN => n5931);
   U1923 : AOI22_X1 port map( A1 => n19410, A2 => n17855, B1 => n19404, B2 => 
                           n18095, ZN => n5909);
   U1924 : AOI22_X1 port map( A1 => n19458, A2 => n17983, B1 => n19452, B2 => 
                           n17759, ZN => n5904);
   U1925 : AOI22_X1 port map( A1 => n19386, A2 => n17713, B1 => n19380, B2 => 
                           n17879, ZN => n5912);
   U1926 : AOI22_X1 port map( A1 => n19187, A2 => n17714, B1 => n19181, B2 => 
                           n17880, ZN => n5867);
   U1927 : AOI22_X1 port map( A1 => n19259, A2 => n17984, B1 => n19253, B2 => 
                           n17760, ZN => n5864);
   U1928 : AOI22_X1 port map( A1 => n19410, A2 => n17856, B1 => n19404, B2 => 
                           n18096, ZN => n5842);
   U1929 : AOI22_X1 port map( A1 => n19458, A2 => n17984, B1 => n19452, B2 => 
                           n17760, ZN => n5837);
   U1930 : AOI22_X1 port map( A1 => n19386, A2 => n17714, B1 => n19380, B2 => 
                           n17880, ZN => n5845);
   U1931 : AOI22_X1 port map( A1 => n19187, A2 => n17715, B1 => n19181, B2 => 
                           n17881, ZN => n5800);
   U1932 : AOI22_X1 port map( A1 => n19259, A2 => n17985, B1 => n19253, B2 => 
                           n17761, ZN => n5797);
   U1933 : AOI22_X1 port map( A1 => n19410, A2 => n17857, B1 => n19404, B2 => 
                           n18097, ZN => n5775);
   U1934 : AOI22_X1 port map( A1 => n19458, A2 => n17985, B1 => n19452, B2 => 
                           n17761, ZN => n5770);
   U1935 : AOI22_X1 port map( A1 => n19386, A2 => n17715, B1 => n19380, B2 => 
                           n17881, ZN => n5778);
   U1936 : AOI22_X1 port map( A1 => n19187, A2 => n17716, B1 => n19181, B2 => 
                           n17882, ZN => n5728);
   U1937 : AOI22_X1 port map( A1 => n19259, A2 => n17986, B1 => n19253, B2 => 
                           n17762, ZN => n5725);
   U1938 : AOI22_X1 port map( A1 => n19410, A2 => n17858, B1 => n19404, B2 => 
                           n18098, ZN => n5703);
   U1939 : AOI22_X1 port map( A1 => n19458, A2 => n17986, B1 => n19452, B2 => 
                           n17762, ZN => n5697);
   U1940 : AOI22_X1 port map( A1 => n19386, A2 => n17716, B1 => n19380, B2 => 
                           n17882, ZN => n5706);
   U1941 : AOI22_X1 port map( A1 => n19187, A2 => n17717, B1 => n19181, B2 => 
                           n17883, ZN => n5658);
   U1942 : AOI22_X1 port map( A1 => n19259, A2 => n17987, B1 => n19253, B2 => 
                           n17763, ZN => n5655);
   U1943 : AOI22_X1 port map( A1 => n19410, A2 => n17859, B1 => n19404, B2 => 
                           n18099, ZN => n5633);
   U1944 : AOI22_X1 port map( A1 => n19458, A2 => n17987, B1 => n19452, B2 => 
                           n17763, ZN => n5626);
   U1945 : AOI22_X1 port map( A1 => n19386, A2 => n17717, B1 => n19380, B2 => 
                           n17883, ZN => n5636);
   U1946 : AOI22_X1 port map( A1 => n19187, A2 => n17718, B1 => n19181, B2 => 
                           n17884, ZN => n5590);
   U1947 : AOI22_X1 port map( A1 => n19259, A2 => n17988, B1 => n19253, B2 => 
                           n17764, ZN => n5587);
   U1948 : AOI22_X1 port map( A1 => n19410, A2 => n17860, B1 => n19404, B2 => 
                           n18100, ZN => n5565);
   U1949 : AOI22_X1 port map( A1 => n19458, A2 => n17988, B1 => n19452, B2 => 
                           n17764, ZN => n5557);
   U1950 : AOI22_X1 port map( A1 => n19386, A2 => n17718, B1 => n19380, B2 => 
                           n17884, ZN => n5568);
   U1951 : AOI22_X1 port map( A1 => n19187, A2 => n17719, B1 => n19181, B2 => 
                           n17885, ZN => n5521);
   U1952 : AOI22_X1 port map( A1 => n19259, A2 => n17989, B1 => n19253, B2 => 
                           n17765, ZN => n5518);
   U1953 : AOI22_X1 port map( A1 => n19410, A2 => n17861, B1 => n19404, B2 => 
                           n18101, ZN => n5496);
   U1954 : AOI22_X1 port map( A1 => n19458, A2 => n17989, B1 => n19452, B2 => 
                           n17765, ZN => n5488);
   U1955 : AOI22_X1 port map( A1 => n19386, A2 => n17719, B1 => n19380, B2 => 
                           n17885, ZN => n5499);
   U1956 : AOI22_X1 port map( A1 => n19187, A2 => n17720, B1 => n19181, B2 => 
                           n17886, ZN => n5452);
   U1957 : AOI22_X1 port map( A1 => n19259, A2 => n17990, B1 => n19253, B2 => 
                           n17766, ZN => n5449);
   U1958 : AOI22_X1 port map( A1 => n19410, A2 => n17862, B1 => n19404, B2 => 
                           n18102, ZN => n5427);
   U1959 : AOI22_X1 port map( A1 => n19458, A2 => n17990, B1 => n19452, B2 => 
                           n17766, ZN => n5420);
   U1960 : AOI22_X1 port map( A1 => n19386, A2 => n17720, B1 => n19380, B2 => 
                           n17886, ZN => n5430);
   U1961 : AOI22_X1 port map( A1 => n19187, A2 => n17721, B1 => n19181, B2 => 
                           n17887, ZN => n5384);
   U1962 : AOI22_X1 port map( A1 => n19259, A2 => n17991, B1 => n19253, B2 => 
                           n17767, ZN => n5381);
   U1963 : AOI22_X1 port map( A1 => n19410, A2 => n17863, B1 => n19404, B2 => 
                           n18103, ZN => n5358);
   U1964 : AOI22_X1 port map( A1 => n19458, A2 => n17991, B1 => n19452, B2 => 
                           n17767, ZN => n5350);
   U1965 : AOI22_X1 port map( A1 => n19386, A2 => n17721, B1 => n19380, B2 => 
                           n17887, ZN => n5362);
   U1966 : AOI22_X1 port map( A1 => n19188, A2 => n17697, B1 => n19182, B2 => 
                           n17912, ZN => n5314);
   U1967 : AOI22_X1 port map( A1 => n19260, A2 => n17992, B1 => n19254, B2 => 
                           n17792, ZN => n5311);
   U1968 : AOI22_X1 port map( A1 => n19459, A2 => n17992, B1 => n19453, B2 => 
                           n17792, ZN => n5121);
   U1969 : AOI22_X1 port map( A1 => n19387, A2 => n17697, B1 => n19381, B2 => 
                           n17912, ZN => n5292);
   U1970 : AOI22_X1 port map( A1 => n19188, A2 => n17698, B1 => n19182, B2 => 
                           n17913, ZN => n4445);
   U1971 : AOI22_X1 port map( A1 => n19260, A2 => n17993, B1 => n19254, B2 => 
                           n17793, ZN => n4378);
   U1972 : AOI22_X1 port map( A1 => n19459, A2 => n17993, B1 => n19453, B2 => 
                           n17793, ZN => n3839);
   U1973 : AOI22_X1 port map( A1 => n19387, A2 => n17698, B1 => n19381, B2 => 
                           n17913, ZN => n4039);
   U1974 : AOI22_X1 port map( A1 => n19188, A2 => n17699, B1 => n19182, B2 => 
                           n17914, ZN => n3286);
   U1975 : AOI22_X1 port map( A1 => n19260, A2 => n17994, B1 => n19254, B2 => 
                           n17794, ZN => n3280);
   U1976 : AOI22_X1 port map( A1 => n19459, A2 => n17994, B1 => n19453, B2 => 
                           n17794, ZN => n3226);
   U1977 : AOI22_X1 port map( A1 => n19387, A2 => n17699, B1 => n19381, B2 => 
                           n17914, ZN => n3242);
   U1978 : AOI22_X1 port map( A1 => n19188, A2 => n17700, B1 => n19182, B2 => 
                           n17915, ZN => n3113);
   U1979 : AOI22_X1 port map( A1 => n19260, A2 => n17995, B1 => n19254, B2 => 
                           n17795, ZN => n3034);
   U1980 : AOI22_X1 port map( A1 => n19459, A2 => n17995, B1 => n19453, B2 => 
                           n17795, ZN => n2782);
   U1981 : AOI22_X1 port map( A1 => n19387, A2 => n17700, B1 => n19381, B2 => 
                           n17915, ZN => n2994);
   U1982 : OAI22_X1 port map( A1 => n19510, A2 => n11487, B1 => n20358, B2 => 
                           n19492, ZN => n7030);
   U1983 : OAI22_X1 port map( A1 => n19510, A2 => n11420, B1 => n20361, B2 => 
                           n19493, ZN => n7034);
   U1984 : OAI22_X1 port map( A1 => n19510, A2 => n11353, B1 => n20364, B2 => 
                           n19494, ZN => n7038);
   U1985 : OAI22_X1 port map( A1 => n19510, A2 => n11286, B1 => n20367, B2 => 
                           n19492, ZN => n7042);
   U1986 : OAI22_X1 port map( A1 => n19509, A2 => n11218, B1 => n20370, B2 => 
                           n19493, ZN => n7046);
   U1987 : OAI22_X1 port map( A1 => n19509, A2 => n11151, B1 => n20373, B2 => 
                           n19494, ZN => n7050);
   U1988 : OAI22_X1 port map( A1 => n19509, A2 => n11084, B1 => n20376, B2 => 
                           n19494, ZN => n7054);
   U1989 : OAI22_X1 port map( A1 => n19509, A2 => n11017, B1 => n20379, B2 => 
                           n19493, ZN => n7058);
   U1990 : OAI22_X1 port map( A1 => n19508, A2 => n10949, B1 => n20382, B2 => 
                           n19494, ZN => n7062);
   U1991 : OAI22_X1 port map( A1 => n19508, A2 => n10882, B1 => n20385, B2 => 
                           n19492, ZN => n7066);
   U1992 : OAI22_X1 port map( A1 => n19508, A2 => n10815, B1 => n20388, B2 => 
                           n19493, ZN => n7070);
   U1993 : OAI22_X1 port map( A1 => n19508, A2 => n10747, B1 => n20391, B2 => 
                           n19492, ZN => n7074);
   U1994 : OAI22_X1 port map( A1 => n19507, A2 => n10680, B1 => n20394, B2 => 
                           n19492, ZN => n7078);
   U1995 : OAI22_X1 port map( A1 => n19507, A2 => n10613, B1 => n20397, B2 => 
                           n19492, ZN => n7082);
   U1996 : OAI22_X1 port map( A1 => n19507, A2 => n10546, B1 => n20400, B2 => 
                           n19492, ZN => n7086);
   U1997 : OAI22_X1 port map( A1 => n19507, A2 => n10478, B1 => n20403, B2 => 
                           n19492, ZN => n7090);
   U1998 : OAI22_X1 port map( A1 => n19506, A2 => n10411, B1 => n20406, B2 => 
                           n19492, ZN => n7094);
   U1999 : OAI22_X1 port map( A1 => n19506, A2 => n10344, B1 => n20409, B2 => 
                           n19492, ZN => n7098);
   U2000 : OAI22_X1 port map( A1 => n19506, A2 => n10277, B1 => n20412, B2 => 
                           n19492, ZN => n7102);
   U2001 : OAI22_X1 port map( A1 => n19506, A2 => n10209, B1 => n20415, B2 => 
                           n19492, ZN => n7106);
   U2002 : OAI22_X1 port map( A1 => n19505, A2 => n10142, B1 => n20418, B2 => 
                           n19492, ZN => n7110);
   U2003 : OAI22_X1 port map( A1 => n19505, A2 => n10075, B1 => n20421, B2 => 
                           n19492, ZN => n7114);
   U2004 : OAI22_X1 port map( A1 => n19505, A2 => n10008, B1 => n20424, B2 => 
                           n19492, ZN => n7118);
   U2005 : OAI22_X1 port map( A1 => n19505, A2 => n9940, B1 => n20427, B2 => 
                           n19493, ZN => n7122);
   U2006 : OAI22_X1 port map( A1 => n19504, A2 => n9873, B1 => n20430, B2 => 
                           n19493, ZN => n7126);
   U2007 : OAI22_X1 port map( A1 => n19504, A2 => n9806, B1 => n20433, B2 => 
                           n19493, ZN => n7130);
   U2008 : OAI22_X1 port map( A1 => n19504, A2 => n9738, B1 => n20436, B2 => 
                           n19493, ZN => n7134);
   U2009 : OAI22_X1 port map( A1 => n19504, A2 => n9671, B1 => n20439, B2 => 
                           n19493, ZN => n7138);
   U2010 : OAI22_X1 port map( A1 => n19503, A2 => n9604, B1 => n20442, B2 => 
                           n19493, ZN => n7142);
   U2011 : OAI22_X1 port map( A1 => n19503, A2 => n9537, B1 => n20445, B2 => 
                           n19493, ZN => n7146);
   U2012 : OAI22_X1 port map( A1 => n19503, A2 => n9469, B1 => n20448, B2 => 
                           n19493, ZN => n7150);
   U2013 : OAI22_X1 port map( A1 => n19502, A2 => n9402, B1 => n20451, B2 => 
                           n19493, ZN => n7154);
   U2014 : OAI22_X1 port map( A1 => n19502, A2 => n9335, B1 => n20454, B2 => 
                           n19493, ZN => n7158);
   U2015 : OAI22_X1 port map( A1 => n19502, A2 => n9268, B1 => n20457, B2 => 
                           n19493, ZN => n7162);
   U2016 : OAI22_X1 port map( A1 => n19502, A2 => n6961, B1 => n20460, B2 => 
                           n19493, ZN => n7166);
   U2017 : OAI22_X1 port map( A1 => n19501, A2 => n6894, B1 => n20463, B2 => 
                           n19493, ZN => n7170);
   U2018 : OAI22_X1 port map( A1 => n19501, A2 => n6827, B1 => n20466, B2 => 
                           n19492, ZN => n7174);
   U2019 : OAI22_X1 port map( A1 => n19501, A2 => n6760, B1 => n20469, B2 => 
                           n19492, ZN => n7178);
   U2020 : OAI22_X1 port map( A1 => n19501, A2 => n6692, B1 => n20472, B2 => 
                           n19494, ZN => n7182);
   U2021 : OAI22_X1 port map( A1 => n19500, A2 => n6625, B1 => n20475, B2 => 
                           n19493, ZN => n7186);
   U2022 : OAI22_X1 port map( A1 => n19500, A2 => n6559, B1 => n20478, B2 => 
                           n19492, ZN => n7190);
   U2023 : OAI22_X1 port map( A1 => n19500, A2 => n6493, B1 => n20481, B2 => 
                           n19492, ZN => n7194);
   U2024 : OAI22_X1 port map( A1 => n19500, A2 => n6427, B1 => n20484, B2 => 
                           n19494, ZN => n7198);
   U2025 : OAI22_X1 port map( A1 => n19499, A2 => n6361, B1 => n20487, B2 => 
                           n19493, ZN => n7202);
   U2026 : OAI22_X1 port map( A1 => n19499, A2 => n6295, B1 => n20490, B2 => 
                           n19492, ZN => n7206);
   U2027 : OAI22_X1 port map( A1 => n19499, A2 => n6229, B1 => n20493, B2 => 
                           n19493, ZN => n7210);
   U2028 : OAI22_X1 port map( A1 => n19499, A2 => n6163, B1 => n20496, B2 => 
                           n19494, ZN => n7214);
   U2029 : OAI22_X1 port map( A1 => n19498, A2 => n6097, B1 => n20499, B2 => 
                           n19494, ZN => n7218);
   U2030 : OAI22_X1 port map( A1 => n19498, A2 => n6029, B1 => n20502, B2 => 
                           n19494, ZN => n7222);
   U2031 : OAI22_X1 port map( A1 => n19498, A2 => n5961, B1 => n20505, B2 => 
                           n19494, ZN => n7226);
   U2032 : OAI22_X1 port map( A1 => n19498, A2 => n5894, B1 => n20508, B2 => 
                           n19494, ZN => n7230);
   U2033 : OAI22_X1 port map( A1 => n19497, A2 => n5827, B1 => n20511, B2 => 
                           n19494, ZN => n7234);
   U2034 : OAI22_X1 port map( A1 => n19497, A2 => n5755, B1 => n20514, B2 => 
                           n19494, ZN => n7238);
   U2035 : OAI22_X1 port map( A1 => n19497, A2 => n5685, B1 => n20517, B2 => 
                           n19494, ZN => n7242);
   U2036 : OAI22_X1 port map( A1 => n19497, A2 => n5617, B1 => n20520, B2 => 
                           n19494, ZN => n7246);
   U2037 : OAI22_X1 port map( A1 => n19496, A2 => n5548, B1 => n20523, B2 => 
                           n19494, ZN => n7250);
   U2038 : OAI22_X1 port map( A1 => n19496, A2 => n5479, B1 => n20526, B2 => 
                           n19494, ZN => n7254);
   U2039 : OAI22_X1 port map( A1 => n19496, A2 => n5411, B1 => n20529, B2 => 
                           n19494, ZN => n7258);
   U2040 : OAI22_X1 port map( A1 => n19495, A2 => n5341, B1 => n20532, B2 => 
                           n19494, ZN => n7262);
   U2041 : INV_X1 port map( A => n2093, ZN => n11716);
   U2042 : OAI22_X1 port map( A1 => n19496, A2 => n4856, B1 => n20535, B2 => 
                           n19493, ZN => n7266);
   U2043 : OAI22_X1 port map( A1 => n19495, A2 => n3638, B1 => n20538, B2 => 
                           n19494, ZN => n7270);
   U2044 : OAI22_X1 port map( A1 => n19495, A2 => n3208, B1 => n20541, B2 => 
                           n19494, ZN => n7274);
   U2045 : OAI22_X1 port map( A1 => n19503, A2 => n2768, B1 => n20572, B2 => 
                           n19492, ZN => n7278);
   U2046 : OAI22_X1 port map( A1 => n20367, A2 => n19578, B1 => n19593, B2 => 
                           n2437, ZN => n7411);
   U2047 : OAI22_X1 port map( A1 => n20370, A2 => n19578, B1 => n19593, B2 => 
                           n2436, ZN => n7412);
   U2048 : OAI22_X1 port map( A1 => n20373, A2 => n19578, B1 => n19593, B2 => 
                           n2435, ZN => n7413);
   U2049 : OAI22_X1 port map( A1 => n20376, A2 => n19578, B1 => n19593, B2 => 
                           n2434, ZN => n7414);
   U2050 : OAI22_X1 port map( A1 => n20379, A2 => n19578, B1 => n19592, B2 => 
                           n2433, ZN => n7415);
   U2051 : OAI22_X1 port map( A1 => n20382, A2 => n19578, B1 => n19592, B2 => 
                           n2432, ZN => n7416);
   U2052 : OAI22_X1 port map( A1 => n20385, A2 => n19578, B1 => n19592, B2 => 
                           n2431, ZN => n7417);
   U2053 : OAI22_X1 port map( A1 => n20388, A2 => n19578, B1 => n19592, B2 => 
                           n2430, ZN => n7418);
   U2054 : OAI22_X1 port map( A1 => n20391, A2 => n19578, B1 => n19591, B2 => 
                           n2429, ZN => n7419);
   U2056 : OAI22_X1 port map( A1 => n20394, A2 => n19578, B1 => n19591, B2 => 
                           n2428, ZN => n7420);
   U2057 : OAI22_X1 port map( A1 => n20397, A2 => n19578, B1 => n19591, B2 => 
                           n2427, ZN => n7421);
   U2058 : OAI22_X1 port map( A1 => n20400, A2 => n19578, B1 => n19591, B2 => 
                           n2426, ZN => n7422);
   U2059 : OAI22_X1 port map( A1 => n20403, A2 => n19577, B1 => n19590, B2 => 
                           n2425, ZN => n7423);
   U2060 : OAI22_X1 port map( A1 => n20406, A2 => n19577, B1 => n19590, B2 => 
                           n2424, ZN => n7424);
   U2061 : OAI22_X1 port map( A1 => n20409, A2 => n19577, B1 => n19590, B2 => 
                           n2423, ZN => n7425);
   U2062 : OAI22_X1 port map( A1 => n20412, A2 => n19577, B1 => n19590, B2 => 
                           n2422, ZN => n7426);
   U2063 : OAI22_X1 port map( A1 => n20415, A2 => n19577, B1 => n19589, B2 => 
                           n2421, ZN => n7427);
   U2064 : OAI22_X1 port map( A1 => n20418, A2 => n19577, B1 => n19589, B2 => 
                           n2420, ZN => n7428);
   U2065 : OAI22_X1 port map( A1 => n20421, A2 => n19577, B1 => n19589, B2 => 
                           n2419, ZN => n7429);
   U2066 : OAI22_X1 port map( A1 => n20424, A2 => n19577, B1 => n19589, B2 => 
                           n2418, ZN => n7430);
   U2067 : OAI22_X1 port map( A1 => n20427, A2 => n19577, B1 => n19588, B2 => 
                           n2417, ZN => n7431);
   U2068 : OAI22_X1 port map( A1 => n20430, A2 => n19577, B1 => n19588, B2 => 
                           n2416, ZN => n7432);
   U2069 : OAI22_X1 port map( A1 => n20433, A2 => n19577, B1 => n19588, B2 => 
                           n2415, ZN => n7433);
   U2070 : OAI22_X1 port map( A1 => n20436, A2 => n19577, B1 => n19588, B2 => 
                           n2414, ZN => n7434);
   U2071 : OAI22_X1 port map( A1 => n20439, A2 => n19576, B1 => n19587, B2 => 
                           n2413, ZN => n7435);
   U2072 : OAI22_X1 port map( A1 => n20442, A2 => n19576, B1 => n19587, B2 => 
                           n2412, ZN => n7436);
   U2073 : OAI22_X1 port map( A1 => n20445, A2 => n19576, B1 => n19587, B2 => 
                           n2411, ZN => n7437);
   U2074 : OAI22_X1 port map( A1 => n20448, A2 => n19576, B1 => n19587, B2 => 
                           n2410, ZN => n7438);
   U2075 : OAI22_X1 port map( A1 => n20451, A2 => n19576, B1 => n19586, B2 => 
                           n2409, ZN => n7439);
   U2076 : OAI22_X1 port map( A1 => n20454, A2 => n19576, B1 => n19586, B2 => 
                           n2408, ZN => n7440);
   U2077 : OAI22_X1 port map( A1 => n20457, A2 => n19576, B1 => n19586, B2 => 
                           n2407, ZN => n7441);
   U2078 : OAI22_X1 port map( A1 => n20460, A2 => n19576, B1 => n19586, B2 => 
                           n2406, ZN => n7442);
   U2079 : OAI22_X1 port map( A1 => n20463, A2 => n19576, B1 => n19585, B2 => 
                           n2405, ZN => n7443);
   U2080 : OAI22_X1 port map( A1 => n20466, A2 => n19576, B1 => n19585, B2 => 
                           n2404, ZN => n7444);
   U2081 : OAI22_X1 port map( A1 => n20469, A2 => n19576, B1 => n19585, B2 => 
                           n2403, ZN => n7445);
   U2082 : OAI22_X1 port map( A1 => n20472, A2 => n19576, B1 => n19585, B2 => 
                           n2402, ZN => n7446);
   U2083 : OAI22_X1 port map( A1 => n20475, A2 => n19578, B1 => n19584, B2 => 
                           n2401, ZN => n7447);
   U2084 : OAI22_X1 port map( A1 => n20478, A2 => n19577, B1 => n19584, B2 => 
                           n2400, ZN => n7448);
   U2085 : OAI22_X1 port map( A1 => n20481, A2 => n19576, B1 => n19584, B2 => 
                           n2399, ZN => n7449);
   U2086 : OAI22_X1 port map( A1 => n20484, A2 => n19578, B1 => n19584, B2 => 
                           n2398, ZN => n7450);
   U2087 : OAI22_X1 port map( A1 => n20487, A2 => n19577, B1 => n19583, B2 => 
                           n2397, ZN => n7451);
   U2088 : OAI22_X1 port map( A1 => n20490, A2 => n19576, B1 => n19583, B2 => 
                           n2396, ZN => n7452);
   U2089 : OAI22_X1 port map( A1 => n20493, A2 => n19578, B1 => n19583, B2 => 
                           n2395, ZN => n7453);
   U2090 : OAI22_X1 port map( A1 => n20496, A2 => n19577, B1 => n19583, B2 => 
                           n2394, ZN => n7454);
   U2091 : OAI22_X1 port map( A1 => n20499, A2 => n19576, B1 => n19582, B2 => 
                           n2393, ZN => n7455);
   U2092 : OAI22_X1 port map( A1 => n20502, A2 => n19578, B1 => n19582, B2 => 
                           n2392, ZN => n7456);
   U2093 : OAI22_X1 port map( A1 => n20505, A2 => n19577, B1 => n19582, B2 => 
                           n2391, ZN => n7457);
   U2094 : OAI22_X1 port map( A1 => n20508, A2 => n19577, B1 => n19582, B2 => 
                           n2390, ZN => n7458);
   U2095 : OAI22_X1 port map( A1 => n20511, A2 => n19578, B1 => n19581, B2 => 
                           n2389, ZN => n7459);
   U2096 : OAI22_X1 port map( A1 => n20514, A2 => n19577, B1 => n19581, B2 => 
                           n2388, ZN => n7460);
   U2097 : OAI22_X1 port map( A1 => n20517, A2 => n19576, B1 => n19581, B2 => 
                           n2387, ZN => n7461);
   U2098 : OAI22_X1 port map( A1 => n20520, A2 => n19576, B1 => n19581, B2 => 
                           n2386, ZN => n7462);
   U2099 : OAI22_X1 port map( A1 => n20523, A2 => n19578, B1 => n19580, B2 => 
                           n2385, ZN => n7463);
   U2100 : OAI22_X1 port map( A1 => n20526, A2 => n19577, B1 => n19580, B2 => 
                           n2384, ZN => n7464);
   U2101 : OAI22_X1 port map( A1 => n20529, A2 => n19576, B1 => n19580, B2 => 
                           n2383, ZN => n7465);
   U2102 : OAI22_X1 port map( A1 => n20532, A2 => n19578, B1 => n19580, B2 => 
                           n2382, ZN => n7466);
   U2103 : OAI22_X1 port map( A1 => n20535, A2 => n19578, B1 => n19579, B2 => 
                           n2381, ZN => n7467);
   U2104 : OAI22_X1 port map( A1 => n20538, A2 => n19577, B1 => n19579, B2 => 
                           n2380, ZN => n7468);
   U2105 : OAI22_X1 port map( A1 => n20541, A2 => n19576, B1 => n19579, B2 => 
                           n2379, ZN => n7469);
   U2106 : OAI22_X1 port map( A1 => n20572, A2 => n19577, B1 => n19579, B2 => 
                           n2378, ZN => n7470);
   U2107 : OAI22_X1 port map( A1 => n20367, A2 => n19802, B1 => n19817, B2 => 
                           n2180, ZN => n7923);
   U2108 : OAI22_X1 port map( A1 => n20370, A2 => n19802, B1 => n19817, B2 => 
                           n2177, ZN => n7924);
   U2109 : OAI22_X1 port map( A1 => n20373, A2 => n19802, B1 => n19817, B2 => 
                           n2174, ZN => n7925);
   U2110 : OAI22_X1 port map( A1 => n20376, A2 => n19802, B1 => n19817, B2 => 
                           n2171, ZN => n7926);
   U2111 : OAI22_X1 port map( A1 => n20379, A2 => n19802, B1 => n19816, B2 => 
                           n2168, ZN => n7927);
   U2112 : OAI22_X1 port map( A1 => n20382, A2 => n19802, B1 => n19816, B2 => 
                           n2165, ZN => n7928);
   U2113 : OAI22_X1 port map( A1 => n20385, A2 => n19802, B1 => n19816, B2 => 
                           n2162, ZN => n7929);
   U2114 : OAI22_X1 port map( A1 => n20388, A2 => n19802, B1 => n19816, B2 => 
                           n2159, ZN => n7930);
   U2115 : OAI22_X1 port map( A1 => n20391, A2 => n19802, B1 => n19815, B2 => 
                           n2156, ZN => n7931);
   U2116 : OAI22_X1 port map( A1 => n20394, A2 => n19802, B1 => n19815, B2 => 
                           n2153, ZN => n7932);
   U2117 : OAI22_X1 port map( A1 => n20397, A2 => n19802, B1 => n19815, B2 => 
                           n2150, ZN => n7933);
   U2118 : OAI22_X1 port map( A1 => n20400, A2 => n19802, B1 => n19815, B2 => 
                           n2147, ZN => n7934);
   U2119 : OAI22_X1 port map( A1 => n20403, A2 => n19801, B1 => n19814, B2 => 
                           n2144, ZN => n7935);
   U2120 : OAI22_X1 port map( A1 => n20406, A2 => n19801, B1 => n19814, B2 => 
                           n2143, ZN => n7936);
   U2121 : OAI22_X1 port map( A1 => n20409, A2 => n19801, B1 => n19814, B2 => 
                           n2142, ZN => n7937);
   U2122 : OAI22_X1 port map( A1 => n20412, A2 => n19801, B1 => n19814, B2 => 
                           n2141, ZN => n7938);
   U2123 : OAI22_X1 port map( A1 => n20415, A2 => n19801, B1 => n19813, B2 => 
                           n2140, ZN => n7939);
   U2124 : OAI22_X1 port map( A1 => n20418, A2 => n19801, B1 => n19813, B2 => 
                           n2139, ZN => n7940);
   U2125 : OAI22_X1 port map( A1 => n20421, A2 => n19801, B1 => n19813, B2 => 
                           n2138, ZN => n7941);
   U2126 : OAI22_X1 port map( A1 => n20424, A2 => n19801, B1 => n19813, B2 => 
                           n2137, ZN => n7942);
   U2127 : OAI22_X1 port map( A1 => n20427, A2 => n19801, B1 => n19812, B2 => 
                           n2136, ZN => n7943);
   U2128 : OAI22_X1 port map( A1 => n20430, A2 => n19801, B1 => n19812, B2 => 
                           n2135, ZN => n7944);
   U2129 : OAI22_X1 port map( A1 => n20433, A2 => n19801, B1 => n19812, B2 => 
                           n2134, ZN => n7945);
   U2130 : OAI22_X1 port map( A1 => n20436, A2 => n19801, B1 => n19812, B2 => 
                           n2133, ZN => n7946);
   U2131 : OAI22_X1 port map( A1 => n20439, A2 => n19800, B1 => n19811, B2 => 
                           n2132, ZN => n7947);
   U2132 : OAI22_X1 port map( A1 => n20442, A2 => n19800, B1 => n19811, B2 => 
                           n2131, ZN => n7948);
   U2133 : OAI22_X1 port map( A1 => n20445, A2 => n19800, B1 => n19811, B2 => 
                           n2130, ZN => n7949);
   U2134 : OAI22_X1 port map( A1 => n20448, A2 => n19800, B1 => n19811, B2 => 
                           n2129, ZN => n7950);
   U2135 : OAI22_X1 port map( A1 => n20451, A2 => n19800, B1 => n19810, B2 => 
                           n2128, ZN => n7951);
   U2136 : OAI22_X1 port map( A1 => n20454, A2 => n19800, B1 => n19810, B2 => 
                           n2127, ZN => n7952);
   U2137 : OAI22_X1 port map( A1 => n20457, A2 => n19800, B1 => n19810, B2 => 
                           n2126, ZN => n7953);
   U2138 : OAI22_X1 port map( A1 => n20460, A2 => n19800, B1 => n19810, B2 => 
                           n2125, ZN => n7954);
   U2139 : OAI22_X1 port map( A1 => n20463, A2 => n19800, B1 => n19809, B2 => 
                           n2124, ZN => n7955);
   U2140 : OAI22_X1 port map( A1 => n20466, A2 => n19800, B1 => n19809, B2 => 
                           n2123, ZN => n7956);
   U2141 : OAI22_X1 port map( A1 => n20469, A2 => n19800, B1 => n19809, B2 => 
                           n2122, ZN => n7957);
   U2142 : OAI22_X1 port map( A1 => n20472, A2 => n19800, B1 => n19809, B2 => 
                           n2121, ZN => n7958);
   U2143 : OAI22_X1 port map( A1 => n20475, A2 => n19802, B1 => n19808, B2 => 
                           n2120, ZN => n7959);
   U2144 : OAI22_X1 port map( A1 => n20478, A2 => n19801, B1 => n19808, B2 => 
                           n2119, ZN => n7960);
   U2145 : OAI22_X1 port map( A1 => n20481, A2 => n19800, B1 => n19808, B2 => 
                           n2118, ZN => n7961);
   U2146 : OAI22_X1 port map( A1 => n20484, A2 => n19802, B1 => n19808, B2 => 
                           n2117, ZN => n7962);
   U2147 : OAI22_X1 port map( A1 => n20487, A2 => n19801, B1 => n19807, B2 => 
                           n2116, ZN => n7963);
   U2148 : OAI22_X1 port map( A1 => n20490, A2 => n19800, B1 => n19807, B2 => 
                           n2115, ZN => n7964);
   U2149 : OAI22_X1 port map( A1 => n20493, A2 => n19802, B1 => n19807, B2 => 
                           n2114, ZN => n7965);
   U2150 : OAI22_X1 port map( A1 => n20496, A2 => n19801, B1 => n19807, B2 => 
                           n2113, ZN => n7966);
   U2151 : OAI22_X1 port map( A1 => n20499, A2 => n19800, B1 => n19806, B2 => 
                           n2112, ZN => n7967);
   U2152 : OAI22_X1 port map( A1 => n20502, A2 => n19802, B1 => n19806, B2 => 
                           n2111, ZN => n7968);
   U2153 : OAI22_X1 port map( A1 => n20505, A2 => n19801, B1 => n19806, B2 => 
                           n2110, ZN => n7969);
   U2154 : OAI22_X1 port map( A1 => n20508, A2 => n19801, B1 => n19806, B2 => 
                           n2109, ZN => n7970);
   U2155 : OAI22_X1 port map( A1 => n20511, A2 => n19802, B1 => n19805, B2 => 
                           n2108, ZN => n7971);
   U2156 : OAI22_X1 port map( A1 => n20514, A2 => n19801, B1 => n19805, B2 => 
                           n2107, ZN => n7972);
   U2157 : OAI22_X1 port map( A1 => n20517, A2 => n19800, B1 => n19805, B2 => 
                           n2106, ZN => n7973);
   U2158 : OAI22_X1 port map( A1 => n20520, A2 => n19800, B1 => n19805, B2 => 
                           n2105, ZN => n7974);
   U2159 : OAI22_X1 port map( A1 => n20523, A2 => n19802, B1 => n19804, B2 => 
                           n2104, ZN => n7975);
   U2160 : OAI22_X1 port map( A1 => n20526, A2 => n19801, B1 => n19804, B2 => 
                           n2103, ZN => n7976);
   U2161 : OAI22_X1 port map( A1 => n20529, A2 => n19800, B1 => n19804, B2 => 
                           n2102, ZN => n7977);
   U2162 : OAI22_X1 port map( A1 => n20532, A2 => n19802, B1 => n19804, B2 => 
                           n2101, ZN => n7978);
   U2163 : OAI22_X1 port map( A1 => n20535, A2 => n19802, B1 => n19803, B2 => 
                           n2100, ZN => n7979);
   U2164 : OAI22_X1 port map( A1 => n20538, A2 => n19801, B1 => n19803, B2 => 
                           n2099, ZN => n7980);
   U2165 : OAI22_X1 port map( A1 => n20541, A2 => n19800, B1 => n19803, B2 => 
                           n2098, ZN => n7981);
   U2166 : OAI22_X1 port map( A1 => n20572, A2 => n19801, B1 => n19803, B2 => 
                           n2097, ZN => n7982);
   U2167 : OAI22_X1 port map( A1 => n20355, A2 => n19493, B1 => n19495, B2 => 
                           n11555, ZN => n7026);
   U2168 : OAI22_X1 port map( A1 => n20368, A2 => n20082, B1 => n20097, B2 => 
                           n1859, ZN => n8563);
   U2169 : OAI22_X1 port map( A1 => n20371, A2 => n20082, B1 => n20097, B2 => 
                           n1858, ZN => n8564);
   U2170 : OAI22_X1 port map( A1 => n20374, A2 => n20082, B1 => n20097, B2 => 
                           n1857, ZN => n8565);
   U2171 : OAI22_X1 port map( A1 => n20377, A2 => n20082, B1 => n20097, B2 => 
                           n1856, ZN => n8566);
   U2172 : OAI22_X1 port map( A1 => n20380, A2 => n20082, B1 => n20096, B2 => 
                           n1855, ZN => n8567);
   U2173 : OAI22_X1 port map( A1 => n20383, A2 => n20082, B1 => n20096, B2 => 
                           n1854, ZN => n8568);
   U2174 : OAI22_X1 port map( A1 => n20386, A2 => n20082, B1 => n20096, B2 => 
                           n1853, ZN => n8569);
   U2175 : OAI22_X1 port map( A1 => n20389, A2 => n20082, B1 => n20096, B2 => 
                           n1852, ZN => n8570);
   U2176 : OAI22_X1 port map( A1 => n20392, A2 => n20082, B1 => n20095, B2 => 
                           n1851, ZN => n8571);
   U2177 : OAI22_X1 port map( A1 => n20395, A2 => n20082, B1 => n20095, B2 => 
                           n1850, ZN => n8572);
   U2178 : OAI22_X1 port map( A1 => n20398, A2 => n20082, B1 => n20095, B2 => 
                           n1849, ZN => n8573);
   U2179 : OAI22_X1 port map( A1 => n20401, A2 => n20082, B1 => n20095, B2 => 
                           n1848, ZN => n8574);
   U2180 : OAI22_X1 port map( A1 => n20404, A2 => n20081, B1 => n20094, B2 => 
                           n1847, ZN => n8575);
   U2181 : OAI22_X1 port map( A1 => n20407, A2 => n20081, B1 => n20094, B2 => 
                           n1846, ZN => n8576);
   U2182 : OAI22_X1 port map( A1 => n20410, A2 => n20081, B1 => n20094, B2 => 
                           n1845, ZN => n8577);
   U2183 : OAI22_X1 port map( A1 => n20413, A2 => n20081, B1 => n20094, B2 => 
                           n1844, ZN => n8578);
   U2184 : OAI22_X1 port map( A1 => n20416, A2 => n20081, B1 => n20093, B2 => 
                           n1843, ZN => n8579);
   U2185 : OAI22_X1 port map( A1 => n20419, A2 => n20081, B1 => n20093, B2 => 
                           n1842, ZN => n8580);
   U2186 : OAI22_X1 port map( A1 => n20422, A2 => n20081, B1 => n20093, B2 => 
                           n1841, ZN => n8581);
   U2187 : OAI22_X1 port map( A1 => n20425, A2 => n20081, B1 => n20093, B2 => 
                           n1840, ZN => n8582);
   U2188 : OAI22_X1 port map( A1 => n20428, A2 => n20081, B1 => n20092, B2 => 
                           n1839, ZN => n8583);
   U2189 : OAI22_X1 port map( A1 => n20431, A2 => n20081, B1 => n20092, B2 => 
                           n1838, ZN => n8584);
   U2190 : OAI22_X1 port map( A1 => n20434, A2 => n20081, B1 => n20092, B2 => 
                           n1837, ZN => n8585);
   U2191 : OAI22_X1 port map( A1 => n20437, A2 => n20081, B1 => n20092, B2 => 
                           n1836, ZN => n8586);
   U2192 : OAI22_X1 port map( A1 => n20440, A2 => n20080, B1 => n20091, B2 => 
                           n1835, ZN => n8587);
   U2193 : OAI22_X1 port map( A1 => n20443, A2 => n20080, B1 => n20091, B2 => 
                           n1834, ZN => n8588);
   U2194 : OAI22_X1 port map( A1 => n20446, A2 => n20080, B1 => n20091, B2 => 
                           n1833, ZN => n8589);
   U2195 : OAI22_X1 port map( A1 => n20449, A2 => n20080, B1 => n20091, B2 => 
                           n1832, ZN => n8590);
   U2196 : OAI22_X1 port map( A1 => n20452, A2 => n20080, B1 => n20090, B2 => 
                           n1831, ZN => n8591);
   U2197 : OAI22_X1 port map( A1 => n20455, A2 => n20080, B1 => n20090, B2 => 
                           n1830, ZN => n8592);
   U2198 : OAI22_X1 port map( A1 => n20458, A2 => n20080, B1 => n20090, B2 => 
                           n1829, ZN => n8593);
   U2199 : OAI22_X1 port map( A1 => n20461, A2 => n20080, B1 => n20090, B2 => 
                           n1828, ZN => n8594);
   U2200 : OAI22_X1 port map( A1 => n20464, A2 => n20080, B1 => n20089, B2 => 
                           n1827, ZN => n8595);
   U2201 : OAI22_X1 port map( A1 => n20467, A2 => n20080, B1 => n20089, B2 => 
                           n1826, ZN => n8596);
   U2202 : OAI22_X1 port map( A1 => n20470, A2 => n20080, B1 => n20089, B2 => 
                           n1825, ZN => n8597);
   U2203 : OAI22_X1 port map( A1 => n20473, A2 => n20080, B1 => n20089, B2 => 
                           n1824, ZN => n8598);
   U2204 : OAI22_X1 port map( A1 => n20476, A2 => n20082, B1 => n20088, B2 => 
                           n1823, ZN => n8599);
   U2205 : OAI22_X1 port map( A1 => n20479, A2 => n20081, B1 => n20088, B2 => 
                           n1822, ZN => n8600);
   U2206 : OAI22_X1 port map( A1 => n20482, A2 => n20080, B1 => n20088, B2 => 
                           n1821, ZN => n8601);
   U2207 : OAI22_X1 port map( A1 => n20485, A2 => n20082, B1 => n20088, B2 => 
                           n1820, ZN => n8602);
   U2208 : OAI22_X1 port map( A1 => n20488, A2 => n20081, B1 => n20087, B2 => 
                           n1819, ZN => n8603);
   U2209 : OAI22_X1 port map( A1 => n20491, A2 => n20080, B1 => n20087, B2 => 
                           n1818, ZN => n8604);
   U2210 : OAI22_X1 port map( A1 => n20494, A2 => n20082, B1 => n20087, B2 => 
                           n1817, ZN => n8605);
   U2211 : OAI22_X1 port map( A1 => n20497, A2 => n20081, B1 => n20087, B2 => 
                           n1816, ZN => n8606);
   U2212 : OAI22_X1 port map( A1 => n20500, A2 => n20080, B1 => n20086, B2 => 
                           n1815, ZN => n8607);
   U2213 : OAI22_X1 port map( A1 => n20503, A2 => n20082, B1 => n20086, B2 => 
                           n1814, ZN => n8608);
   U2214 : OAI22_X1 port map( A1 => n20506, A2 => n20081, B1 => n20086, B2 => 
                           n1813, ZN => n8609);
   U2215 : OAI22_X1 port map( A1 => n20509, A2 => n20081, B1 => n20086, B2 => 
                           n1812, ZN => n8610);
   U2216 : OAI22_X1 port map( A1 => n20512, A2 => n20082, B1 => n20085, B2 => 
                           n1811, ZN => n8611);
   U2217 : OAI22_X1 port map( A1 => n20515, A2 => n20081, B1 => n20085, B2 => 
                           n1810, ZN => n8612);
   U2218 : OAI22_X1 port map( A1 => n20518, A2 => n20080, B1 => n20085, B2 => 
                           n1809, ZN => n8613);
   U2219 : OAI22_X1 port map( A1 => n20521, A2 => n20080, B1 => n20085, B2 => 
                           n1808, ZN => n8614);
   U2220 : OAI22_X1 port map( A1 => n20524, A2 => n20082, B1 => n20084, B2 => 
                           n1807, ZN => n8615);
   U2221 : OAI22_X1 port map( A1 => n20527, A2 => n20081, B1 => n20084, B2 => 
                           n1806, ZN => n8616);
   U2222 : OAI22_X1 port map( A1 => n20530, A2 => n20080, B1 => n20084, B2 => 
                           n1805, ZN => n8617);
   U2223 : OAI22_X1 port map( A1 => n20533, A2 => n20082, B1 => n20084, B2 => 
                           n1804, ZN => n8618);
   U2224 : OAI22_X1 port map( A1 => n20536, A2 => n20082, B1 => n20083, B2 => 
                           n1803, ZN => n8619);
   U2225 : OAI22_X1 port map( A1 => n20539, A2 => n20081, B1 => n20083, B2 => 
                           n1802, ZN => n8620);
   U2226 : OAI22_X1 port map( A1 => n20542, A2 => n20080, B1 => n20083, B2 => 
                           n1801, ZN => n8621);
   U2227 : OAI22_X1 port map( A1 => n20573, A2 => n20081, B1 => n20083, B2 => 
                           n1800, ZN => n8622);
   U2228 : OAI22_X1 port map( A1 => n20368, A2 => n20110, B1 => n20125, B2 => 
                           n1792, ZN => n8627);
   U2229 : OAI22_X1 port map( A1 => n20371, A2 => n20110, B1 => n20125, B2 => 
                           n1791, ZN => n8628);
   U2230 : OAI22_X1 port map( A1 => n20374, A2 => n20110, B1 => n20125, B2 => 
                           n1790, ZN => n8629);
   U2231 : OAI22_X1 port map( A1 => n20377, A2 => n20110, B1 => n20125, B2 => 
                           n1789, ZN => n8630);
   U2232 : OAI22_X1 port map( A1 => n20380, A2 => n20110, B1 => n20124, B2 => 
                           n1788, ZN => n8631);
   U2233 : OAI22_X1 port map( A1 => n20383, A2 => n20110, B1 => n20124, B2 => 
                           n1787, ZN => n8632);
   U2234 : OAI22_X1 port map( A1 => n20386, A2 => n20110, B1 => n20124, B2 => 
                           n1786, ZN => n8633);
   U2235 : OAI22_X1 port map( A1 => n20389, A2 => n20110, B1 => n20124, B2 => 
                           n1785, ZN => n8634);
   U2236 : OAI22_X1 port map( A1 => n20392, A2 => n20110, B1 => n20123, B2 => 
                           n1784, ZN => n8635);
   U2237 : OAI22_X1 port map( A1 => n20395, A2 => n20110, B1 => n20123, B2 => 
                           n1783, ZN => n8636);
   U2238 : OAI22_X1 port map( A1 => n20398, A2 => n20110, B1 => n20123, B2 => 
                           n1782, ZN => n8637);
   U2239 : OAI22_X1 port map( A1 => n20401, A2 => n20110, B1 => n20123, B2 => 
                           n1781, ZN => n8638);
   U2240 : OAI22_X1 port map( A1 => n20404, A2 => n20109, B1 => n20122, B2 => 
                           n1780, ZN => n8639);
   U2241 : OAI22_X1 port map( A1 => n20407, A2 => n20109, B1 => n20122, B2 => 
                           n1779, ZN => n8640);
   U2242 : OAI22_X1 port map( A1 => n20410, A2 => n20109, B1 => n20122, B2 => 
                           n1778, ZN => n8641);
   U2243 : OAI22_X1 port map( A1 => n20413, A2 => n20109, B1 => n20122, B2 => 
                           n1777, ZN => n8642);
   U2244 : OAI22_X1 port map( A1 => n20416, A2 => n20109, B1 => n20121, B2 => 
                           n1776, ZN => n8643);
   U2245 : OAI22_X1 port map( A1 => n20419, A2 => n20109, B1 => n20121, B2 => 
                           n1775, ZN => n8644);
   U2246 : OAI22_X1 port map( A1 => n20422, A2 => n20109, B1 => n20121, B2 => 
                           n1774, ZN => n8645);
   U2247 : OAI22_X1 port map( A1 => n20425, A2 => n20109, B1 => n20121, B2 => 
                           n1773, ZN => n8646);
   U2248 : OAI22_X1 port map( A1 => n20428, A2 => n20109, B1 => n20120, B2 => 
                           n1772, ZN => n8647);
   U2249 : OAI22_X1 port map( A1 => n20431, A2 => n20109, B1 => n20120, B2 => 
                           n1771, ZN => n8648);
   U2250 : OAI22_X1 port map( A1 => n20434, A2 => n20109, B1 => n20120, B2 => 
                           n1770, ZN => n8649);
   U2251 : OAI22_X1 port map( A1 => n20437, A2 => n20109, B1 => n20120, B2 => 
                           n1769, ZN => n8650);
   U2252 : OAI22_X1 port map( A1 => n20440, A2 => n20108, B1 => n20119, B2 => 
                           n1768, ZN => n8651);
   U2253 : OAI22_X1 port map( A1 => n20443, A2 => n20108, B1 => n20119, B2 => 
                           n1767, ZN => n8652);
   U2254 : OAI22_X1 port map( A1 => n20446, A2 => n20108, B1 => n20119, B2 => 
                           n1766, ZN => n8653);
   U2255 : OAI22_X1 port map( A1 => n20449, A2 => n20108, B1 => n20119, B2 => 
                           n1765, ZN => n8654);
   U2256 : OAI22_X1 port map( A1 => n20452, A2 => n20108, B1 => n20118, B2 => 
                           n1764, ZN => n8655);
   U2257 : OAI22_X1 port map( A1 => n20455, A2 => n20108, B1 => n20118, B2 => 
                           n1763, ZN => n8656);
   U2258 : OAI22_X1 port map( A1 => n20458, A2 => n20108, B1 => n20118, B2 => 
                           n1762, ZN => n8657);
   U2259 : OAI22_X1 port map( A1 => n20461, A2 => n20108, B1 => n20118, B2 => 
                           n1761, ZN => n8658);
   U2260 : OAI22_X1 port map( A1 => n20464, A2 => n20108, B1 => n20117, B2 => 
                           n1760, ZN => n8659);
   U2261 : OAI22_X1 port map( A1 => n20467, A2 => n20108, B1 => n20117, B2 => 
                           n1759, ZN => n8660);
   U2262 : OAI22_X1 port map( A1 => n20470, A2 => n20108, B1 => n20117, B2 => 
                           n1758, ZN => n8661);
   U2263 : OAI22_X1 port map( A1 => n20473, A2 => n20108, B1 => n20117, B2 => 
                           n1757, ZN => n8662);
   U2264 : OAI22_X1 port map( A1 => n20476, A2 => n20110, B1 => n20116, B2 => 
                           n1756, ZN => n8663);
   U2265 : OAI22_X1 port map( A1 => n20479, A2 => n20109, B1 => n20116, B2 => 
                           n1755, ZN => n8664);
   U2266 : OAI22_X1 port map( A1 => n20482, A2 => n20108, B1 => n20116, B2 => 
                           n1754, ZN => n8665);
   U2267 : OAI22_X1 port map( A1 => n20485, A2 => n20110, B1 => n20116, B2 => 
                           n1753, ZN => n8666);
   U2268 : OAI22_X1 port map( A1 => n20488, A2 => n20109, B1 => n20115, B2 => 
                           n1752, ZN => n8667);
   U2269 : OAI22_X1 port map( A1 => n20491, A2 => n20108, B1 => n20115, B2 => 
                           n1751, ZN => n8668);
   U2270 : OAI22_X1 port map( A1 => n20494, A2 => n20110, B1 => n20115, B2 => 
                           n1750, ZN => n8669);
   U2271 : OAI22_X1 port map( A1 => n20497, A2 => n20109, B1 => n20115, B2 => 
                           n1749, ZN => n8670);
   U2272 : OAI22_X1 port map( A1 => n20500, A2 => n20108, B1 => n20114, B2 => 
                           n1745, ZN => n8671);
   U2273 : OAI22_X1 port map( A1 => n20503, A2 => n20110, B1 => n20114, B2 => 
                           n1744, ZN => n8672);
   U2274 : OAI22_X1 port map( A1 => n20506, A2 => n20109, B1 => n20114, B2 => 
                           n1743, ZN => n8673);
   U2275 : OAI22_X1 port map( A1 => n20509, A2 => n20109, B1 => n20114, B2 => 
                           n1742, ZN => n8674);
   U2276 : OAI22_X1 port map( A1 => n20512, A2 => n20110, B1 => n20113, B2 => 
                           n1741, ZN => n8675);
   U2277 : OAI22_X1 port map( A1 => n20515, A2 => n20109, B1 => n20113, B2 => 
                           n1740, ZN => n8676);
   U2278 : OAI22_X1 port map( A1 => n20518, A2 => n20108, B1 => n20113, B2 => 
                           n1739, ZN => n8677);
   U2279 : OAI22_X1 port map( A1 => n20521, A2 => n20108, B1 => n20113, B2 => 
                           n1738, ZN => n8678);
   U2280 : OAI22_X1 port map( A1 => n20524, A2 => n20110, B1 => n20112, B2 => 
                           n1737, ZN => n8679);
   U2281 : OAI22_X1 port map( A1 => n20527, A2 => n20109, B1 => n20112, B2 => 
                           n1736, ZN => n8680);
   U2282 : OAI22_X1 port map( A1 => n20530, A2 => n20108, B1 => n20112, B2 => 
                           n1735, ZN => n8681);
   U2283 : OAI22_X1 port map( A1 => n20533, A2 => n20110, B1 => n20112, B2 => 
                           n1734, ZN => n8682);
   U2284 : OAI22_X1 port map( A1 => n20536, A2 => n20110, B1 => n20111, B2 => 
                           n1733, ZN => n8683);
   U2285 : OAI22_X1 port map( A1 => n20539, A2 => n20109, B1 => n20111, B2 => 
                           n1732, ZN => n8684);
   U2286 : OAI22_X1 port map( A1 => n20542, A2 => n20108, B1 => n20111, B2 => 
                           n1731, ZN => n8685);
   U2287 : OAI22_X1 port map( A1 => n20573, A2 => n20109, B1 => n20111, B2 => 
                           n1730, ZN => n8686);
   U2288 : OAI22_X1 port map( A1 => n20355, A2 => n19577, B1 => n19594, B2 => 
                           n2441, ZN => n7407);
   U2289 : OAI22_X1 port map( A1 => n20358, A2 => n19576, B1 => n19594, B2 => 
                           n2440, ZN => n7408);
   U2290 : OAI22_X1 port map( A1 => n20361, A2 => n19576, B1 => n19594, B2 => 
                           n2439, ZN => n7409);
   U2291 : OAI22_X1 port map( A1 => n20364, A2 => n19578, B1 => n19594, B2 => 
                           n2438, ZN => n7410);
   U2292 : OAI22_X1 port map( A1 => n20355, A2 => n19801, B1 => n19818, B2 => 
                           n2192, ZN => n7919);
   U2293 : OAI22_X1 port map( A1 => n20358, A2 => n19800, B1 => n19818, B2 => 
                           n2189, ZN => n7920);
   U2294 : OAI22_X1 port map( A1 => n20361, A2 => n19800, B1 => n19818, B2 => 
                           n2186, ZN => n7921);
   U2295 : OAI22_X1 port map( A1 => n20364, A2 => n19802, B1 => n19818, B2 => 
                           n2183, ZN => n7922);
   U2296 : OAI22_X1 port map( A1 => n20356, A2 => n20081, B1 => n20098, B2 => 
                           n1863, ZN => n8559);
   U2297 : OAI22_X1 port map( A1 => n20359, A2 => n20080, B1 => n20098, B2 => 
                           n1862, ZN => n8560);
   U2298 : OAI22_X1 port map( A1 => n20362, A2 => n20080, B1 => n20098, B2 => 
                           n1861, ZN => n8561);
   U2299 : OAI22_X1 port map( A1 => n20365, A2 => n20082, B1 => n20098, B2 => 
                           n1860, ZN => n8562);
   U2300 : OAI22_X1 port map( A1 => n20356, A2 => n20109, B1 => n20126, B2 => 
                           n1796, ZN => n8623);
   U2301 : OAI22_X1 port map( A1 => n20359, A2 => n20108, B1 => n20126, B2 => 
                           n1795, ZN => n8624);
   U2302 : OAI22_X1 port map( A1 => n20362, A2 => n20108, B1 => n20126, B2 => 
                           n1794, ZN => n8625);
   U2303 : OAI22_X1 port map( A1 => n20365, A2 => n20110, B1 => n20126, B2 => 
                           n1793, ZN => n8626);
   U2304 : OAI22_X1 port map( A1 => n20367, A2 => n19550, B1 => n19565, B2 => 
                           n2759, ZN => n7347);
   U2305 : OAI22_X1 port map( A1 => n20370, A2 => n19550, B1 => n19565, B2 => 
                           n2758, ZN => n7348);
   U2306 : OAI22_X1 port map( A1 => n20373, A2 => n19550, B1 => n19565, B2 => 
                           n2757, ZN => n7349);
   U2307 : OAI22_X1 port map( A1 => n20376, A2 => n19550, B1 => n19565, B2 => 
                           n2756, ZN => n7350);
   U2308 : OAI22_X1 port map( A1 => n20379, A2 => n19550, B1 => n19564, B2 => 
                           n2755, ZN => n7351);
   U2309 : OAI22_X1 port map( A1 => n20382, A2 => n19550, B1 => n19564, B2 => 
                           n2754, ZN => n7352);
   U2310 : OAI22_X1 port map( A1 => n20385, A2 => n19550, B1 => n19564, B2 => 
                           n2753, ZN => n7353);
   U2311 : OAI22_X1 port map( A1 => n20388, A2 => n19550, B1 => n19564, B2 => 
                           n2752, ZN => n7354);
   U2312 : OAI22_X1 port map( A1 => n20391, A2 => n19550, B1 => n19563, B2 => 
                           n2751, ZN => n7355);
   U2313 : OAI22_X1 port map( A1 => n20394, A2 => n19550, B1 => n19563, B2 => 
                           n2750, ZN => n7356);
   U2314 : OAI22_X1 port map( A1 => n20397, A2 => n19550, B1 => n19563, B2 => 
                           n2749, ZN => n7357);
   U2315 : OAI22_X1 port map( A1 => n20400, A2 => n19550, B1 => n19563, B2 => 
                           n2748, ZN => n7358);
   U2316 : OAI22_X1 port map( A1 => n20403, A2 => n19549, B1 => n19562, B2 => 
                           n2747, ZN => n7359);
   U2317 : OAI22_X1 port map( A1 => n20406, A2 => n19549, B1 => n19562, B2 => 
                           n2746, ZN => n7360);
   U2318 : OAI22_X1 port map( A1 => n20409, A2 => n19549, B1 => n19562, B2 => 
                           n2745, ZN => n7361);
   U2319 : OAI22_X1 port map( A1 => n20412, A2 => n19549, B1 => n19562, B2 => 
                           n2744, ZN => n7362);
   U2320 : OAI22_X1 port map( A1 => n20415, A2 => n19549, B1 => n19561, B2 => 
                           n2743, ZN => n7363);
   U2321 : OAI22_X1 port map( A1 => n20418, A2 => n19549, B1 => n19561, B2 => 
                           n2742, ZN => n7364);
   U2322 : OAI22_X1 port map( A1 => n20421, A2 => n19549, B1 => n19561, B2 => 
                           n2741, ZN => n7365);
   U2323 : OAI22_X1 port map( A1 => n20424, A2 => n19549, B1 => n19561, B2 => 
                           n2740, ZN => n7366);
   U2324 : OAI22_X1 port map( A1 => n20427, A2 => n19549, B1 => n19560, B2 => 
                           n2739, ZN => n7367);
   U2325 : OAI22_X1 port map( A1 => n20430, A2 => n19549, B1 => n19560, B2 => 
                           n2738, ZN => n7368);
   U2326 : OAI22_X1 port map( A1 => n20433, A2 => n19549, B1 => n19560, B2 => 
                           n2737, ZN => n7369);
   U2327 : OAI22_X1 port map( A1 => n20436, A2 => n19549, B1 => n19560, B2 => 
                           n2736, ZN => n7370);
   U2328 : OAI22_X1 port map( A1 => n20439, A2 => n19548, B1 => n19559, B2 => 
                           n2735, ZN => n7371);
   U2329 : OAI22_X1 port map( A1 => n20442, A2 => n19548, B1 => n19559, B2 => 
                           n2734, ZN => n7372);
   U2330 : OAI22_X1 port map( A1 => n20445, A2 => n19548, B1 => n19559, B2 => 
                           n2733, ZN => n7373);
   U2331 : OAI22_X1 port map( A1 => n20448, A2 => n19548, B1 => n19559, B2 => 
                           n2732, ZN => n7374);
   U2332 : OAI22_X1 port map( A1 => n20451, A2 => n19548, B1 => n19558, B2 => 
                           n2731, ZN => n7375);
   U2333 : OAI22_X1 port map( A1 => n20454, A2 => n19548, B1 => n19558, B2 => 
                           n2730, ZN => n7376);
   U2334 : OAI22_X1 port map( A1 => n20457, A2 => n19548, B1 => n19558, B2 => 
                           n2729, ZN => n7377);
   U2335 : OAI22_X1 port map( A1 => n20460, A2 => n19548, B1 => n19558, B2 => 
                           n2728, ZN => n7378);
   U2336 : OAI22_X1 port map( A1 => n20463, A2 => n19548, B1 => n19557, B2 => 
                           n2727, ZN => n7379);
   U2337 : OAI22_X1 port map( A1 => n20466, A2 => n19548, B1 => n19557, B2 => 
                           n2726, ZN => n7380);
   U2338 : OAI22_X1 port map( A1 => n20469, A2 => n19548, B1 => n19557, B2 => 
                           n2725, ZN => n7381);
   U2339 : OAI22_X1 port map( A1 => n20472, A2 => n19548, B1 => n19557, B2 => 
                           n2724, ZN => n7382);
   U2340 : OAI22_X1 port map( A1 => n20475, A2 => n19550, B1 => n19556, B2 => 
                           n2723, ZN => n7383);
   U2341 : OAI22_X1 port map( A1 => n20478, A2 => n19549, B1 => n19556, B2 => 
                           n2722, ZN => n7384);
   U2342 : OAI22_X1 port map( A1 => n20481, A2 => n19548, B1 => n19556, B2 => 
                           n2721, ZN => n7385);
   U2343 : OAI22_X1 port map( A1 => n20484, A2 => n19550, B1 => n19556, B2 => 
                           n2720, ZN => n7386);
   U2344 : OAI22_X1 port map( A1 => n20487, A2 => n19549, B1 => n19555, B2 => 
                           n2463, ZN => n7387);
   U2345 : OAI22_X1 port map( A1 => n20490, A2 => n19548, B1 => n19555, B2 => 
                           n2462, ZN => n7388);
   U2346 : OAI22_X1 port map( A1 => n20493, A2 => n19550, B1 => n19555, B2 => 
                           n2461, ZN => n7389);
   U2347 : OAI22_X1 port map( A1 => n20496, A2 => n19549, B1 => n19555, B2 => 
                           n2460, ZN => n7390);
   U2348 : OAI22_X1 port map( A1 => n20499, A2 => n19548, B1 => n19554, B2 => 
                           n2459, ZN => n7391);
   U2349 : OAI22_X1 port map( A1 => n20502, A2 => n19550, B1 => n19554, B2 => 
                           n2458, ZN => n7392);
   U2350 : OAI22_X1 port map( A1 => n20505, A2 => n19549, B1 => n19554, B2 => 
                           n2457, ZN => n7393);
   U2351 : OAI22_X1 port map( A1 => n20508, A2 => n19549, B1 => n19554, B2 => 
                           n2456, ZN => n7394);
   U2352 : OAI22_X1 port map( A1 => n20511, A2 => n19550, B1 => n19553, B2 => 
                           n2455, ZN => n7395);
   U2353 : OAI22_X1 port map( A1 => n20514, A2 => n19549, B1 => n19553, B2 => 
                           n2454, ZN => n7396);
   U2354 : OAI22_X1 port map( A1 => n20517, A2 => n19548, B1 => n19553, B2 => 
                           n2453, ZN => n7397);
   U2355 : OAI22_X1 port map( A1 => n20520, A2 => n19548, B1 => n19553, B2 => 
                           n2452, ZN => n7398);
   U2356 : OAI22_X1 port map( A1 => n20523, A2 => n19550, B1 => n19552, B2 => 
                           n2451, ZN => n7399);
   U2357 : OAI22_X1 port map( A1 => n20526, A2 => n19549, B1 => n19552, B2 => 
                           n2450, ZN => n7400);
   U2358 : OAI22_X1 port map( A1 => n20529, A2 => n19548, B1 => n19552, B2 => 
                           n2449, ZN => n7401);
   U2359 : OAI22_X1 port map( A1 => n20532, A2 => n19550, B1 => n19552, B2 => 
                           n2448, ZN => n7402);
   U2360 : OAI22_X1 port map( A1 => n20535, A2 => n19550, B1 => n19551, B2 => 
                           n2447, ZN => n7403);
   U2361 : OAI22_X1 port map( A1 => n20538, A2 => n19549, B1 => n19551, B2 => 
                           n2446, ZN => n7404);
   U2362 : OAI22_X1 port map( A1 => n20541, A2 => n19548, B1 => n19551, B2 => 
                           n2445, ZN => n7405);
   U2363 : OAI22_X1 port map( A1 => n20572, A2 => n19549, B1 => n19551, B2 => 
                           n2444, ZN => n7406);
   U2364 : OAI22_X1 port map( A1 => n20368, A2 => n19998, B1 => n20013, B2 => 
                           n1933, ZN => n8371);
   U2365 : OAI22_X1 port map( A1 => n20371, A2 => n19998, B1 => n20013, B2 => 
                           n1932, ZN => n8372);
   U2366 : OAI22_X1 port map( A1 => n20374, A2 => n19998, B1 => n20013, B2 => 
                           n1931, ZN => n8373);
   U2367 : OAI22_X1 port map( A1 => n20377, A2 => n19998, B1 => n20013, B2 => 
                           n1930, ZN => n8374);
   U2368 : OAI22_X1 port map( A1 => n20380, A2 => n19998, B1 => n20012, B2 => 
                           n1929, ZN => n8375);
   U2369 : OAI22_X1 port map( A1 => n20383, A2 => n19998, B1 => n20012, B2 => 
                           n1928, ZN => n8376);
   U2370 : OAI22_X1 port map( A1 => n20386, A2 => n19998, B1 => n20012, B2 => 
                           n1927, ZN => n8377);
   U2371 : OAI22_X1 port map( A1 => n20389, A2 => n19998, B1 => n20012, B2 => 
                           n1926, ZN => n8378);
   U2372 : OAI22_X1 port map( A1 => n20392, A2 => n19998, B1 => n20011, B2 => 
                           n1925, ZN => n8379);
   U2373 : OAI22_X1 port map( A1 => n20395, A2 => n19998, B1 => n20011, B2 => 
                           n1924, ZN => n8380);
   U2374 : OAI22_X1 port map( A1 => n20398, A2 => n19998, B1 => n20011, B2 => 
                           n1923, ZN => n8381);
   U2375 : OAI22_X1 port map( A1 => n20401, A2 => n19998, B1 => n20011, B2 => 
                           n1922, ZN => n8382);
   U2376 : OAI22_X1 port map( A1 => n20404, A2 => n19997, B1 => n20010, B2 => 
                           n1921, ZN => n8383);
   U2377 : OAI22_X1 port map( A1 => n20407, A2 => n19997, B1 => n20010, B2 => 
                           n1920, ZN => n8384);
   U2378 : OAI22_X1 port map( A1 => n20410, A2 => n19997, B1 => n20010, B2 => 
                           n1919, ZN => n8385);
   U2379 : OAI22_X1 port map( A1 => n20413, A2 => n19997, B1 => n20010, B2 => 
                           n1918, ZN => n8386);
   U2380 : OAI22_X1 port map( A1 => n20416, A2 => n19997, B1 => n20009, B2 => 
                           n1917, ZN => n8387);
   U2381 : OAI22_X1 port map( A1 => n20419, A2 => n19997, B1 => n20009, B2 => 
                           n1916, ZN => n8388);
   U2382 : OAI22_X1 port map( A1 => n20422, A2 => n19997, B1 => n20009, B2 => 
                           n1915, ZN => n8389);
   U2383 : OAI22_X1 port map( A1 => n20425, A2 => n19997, B1 => n20009, B2 => 
                           n1914, ZN => n8390);
   U2384 : OAI22_X1 port map( A1 => n20428, A2 => n19997, B1 => n20008, B2 => 
                           n1913, ZN => n8391);
   U2385 : OAI22_X1 port map( A1 => n20431, A2 => n19997, B1 => n20008, B2 => 
                           n1912, ZN => n8392);
   U2386 : OAI22_X1 port map( A1 => n20434, A2 => n19997, B1 => n20008, B2 => 
                           n1911, ZN => n8393);
   U2387 : OAI22_X1 port map( A1 => n20437, A2 => n19997, B1 => n20008, B2 => 
                           n1910, ZN => n8394);
   U2388 : OAI22_X1 port map( A1 => n20440, A2 => n19996, B1 => n20007, B2 => 
                           n1909, ZN => n8395);
   U2389 : OAI22_X1 port map( A1 => n20443, A2 => n19996, B1 => n20007, B2 => 
                           n1908, ZN => n8396);
   U2390 : OAI22_X1 port map( A1 => n20446, A2 => n19996, B1 => n20007, B2 => 
                           n1907, ZN => n8397);
   U2391 : OAI22_X1 port map( A1 => n20449, A2 => n19996, B1 => n20007, B2 => 
                           n1906, ZN => n8398);
   U2392 : OAI22_X1 port map( A1 => n20452, A2 => n19996, B1 => n20006, B2 => 
                           n1905, ZN => n8399);
   U2393 : OAI22_X1 port map( A1 => n20455, A2 => n19996, B1 => n20006, B2 => 
                           n1904, ZN => n8400);
   U2394 : OAI22_X1 port map( A1 => n20458, A2 => n19996, B1 => n20006, B2 => 
                           n1903, ZN => n8401);
   U2395 : OAI22_X1 port map( A1 => n20461, A2 => n19996, B1 => n20006, B2 => 
                           n1902, ZN => n8402);
   U2396 : OAI22_X1 port map( A1 => n20464, A2 => n19996, B1 => n20005, B2 => 
                           n1901, ZN => n8403);
   U2397 : OAI22_X1 port map( A1 => n20467, A2 => n19996, B1 => n20005, B2 => 
                           n1900, ZN => n8404);
   U2398 : OAI22_X1 port map( A1 => n20470, A2 => n19996, B1 => n20005, B2 => 
                           n1899, ZN => n8405);
   U2399 : OAI22_X1 port map( A1 => n20473, A2 => n19996, B1 => n20005, B2 => 
                           n1898, ZN => n8406);
   U2400 : OAI22_X1 port map( A1 => n20476, A2 => n19998, B1 => n20004, B2 => 
                           n1897, ZN => n8407);
   U2401 : OAI22_X1 port map( A1 => n20479, A2 => n19997, B1 => n20004, B2 => 
                           n1896, ZN => n8408);
   U2402 : OAI22_X1 port map( A1 => n20482, A2 => n19996, B1 => n20004, B2 => 
                           n1895, ZN => n8409);
   U2403 : OAI22_X1 port map( A1 => n20485, A2 => n19998, B1 => n20004, B2 => 
                           n1894, ZN => n8410);
   U2404 : OAI22_X1 port map( A1 => n20488, A2 => n19997, B1 => n20003, B2 => 
                           n1893, ZN => n8411);
   U2405 : OAI22_X1 port map( A1 => n20491, A2 => n19996, B1 => n20003, B2 => 
                           n1892, ZN => n8412);
   U2406 : OAI22_X1 port map( A1 => n20494, A2 => n19998, B1 => n20003, B2 => 
                           n1891, ZN => n8413);
   U2407 : OAI22_X1 port map( A1 => n20497, A2 => n19997, B1 => n20003, B2 => 
                           n1890, ZN => n8414);
   U2408 : OAI22_X1 port map( A1 => n20500, A2 => n19996, B1 => n20002, B2 => 
                           n1889, ZN => n8415);
   U2409 : OAI22_X1 port map( A1 => n20503, A2 => n19998, B1 => n20002, B2 => 
                           n1888, ZN => n8416);
   U2410 : OAI22_X1 port map( A1 => n20506, A2 => n19997, B1 => n20002, B2 => 
                           n1887, ZN => n8417);
   U2411 : OAI22_X1 port map( A1 => n20509, A2 => n19997, B1 => n20002, B2 => 
                           n1886, ZN => n8418);
   U2412 : OAI22_X1 port map( A1 => n20512, A2 => n19998, B1 => n20001, B2 => 
                           n1885, ZN => n8419);
   U2413 : OAI22_X1 port map( A1 => n20515, A2 => n19997, B1 => n20001, B2 => 
                           n1884, ZN => n8420);
   U2414 : OAI22_X1 port map( A1 => n20518, A2 => n19996, B1 => n20001, B2 => 
                           n1883, ZN => n8421);
   U2415 : OAI22_X1 port map( A1 => n20521, A2 => n19996, B1 => n20001, B2 => 
                           n1882, ZN => n8422);
   U2416 : OAI22_X1 port map( A1 => n20524, A2 => n19998, B1 => n20000, B2 => 
                           n1881, ZN => n8423);
   U2417 : OAI22_X1 port map( A1 => n20527, A2 => n19997, B1 => n20000, B2 => 
                           n1880, ZN => n8424);
   U2418 : OAI22_X1 port map( A1 => n20530, A2 => n19996, B1 => n20000, B2 => 
                           n1879, ZN => n8425);
   U2419 : OAI22_X1 port map( A1 => n20533, A2 => n19998, B1 => n20000, B2 => 
                           n1878, ZN => n8426);
   U2420 : OAI22_X1 port map( A1 => n20536, A2 => n19998, B1 => n19999, B2 => 
                           n1877, ZN => n8427);
   U2421 : OAI22_X1 port map( A1 => n20539, A2 => n19997, B1 => n19999, B2 => 
                           n1876, ZN => n8428);
   U2422 : OAI22_X1 port map( A1 => n20542, A2 => n19996, B1 => n19999, B2 => 
                           n1875, ZN => n8429);
   U2423 : OAI22_X1 port map( A1 => n20573, A2 => n19997, B1 => n19999, B2 => 
                           n1874, ZN => n8430);
   U2424 : OAI22_X1 port map( A1 => n20355, A2 => n19549, B1 => n19566, B2 => 
                           n2763, ZN => n7343);
   U2425 : OAI22_X1 port map( A1 => n20358, A2 => n19548, B1 => n19566, B2 => 
                           n2762, ZN => n7344);
   U2426 : OAI22_X1 port map( A1 => n20361, A2 => n19548, B1 => n19566, B2 => 
                           n2761, ZN => n7345);
   U2427 : OAI22_X1 port map( A1 => n20364, A2 => n19550, B1 => n19566, B2 => 
                           n2760, ZN => n7346);
   U2428 : OAI22_X1 port map( A1 => n20356, A2 => n19997, B1 => n20014, B2 => 
                           n1937, ZN => n8367);
   U2429 : OAI22_X1 port map( A1 => n20359, A2 => n19996, B1 => n20014, B2 => 
                           n1936, ZN => n8368);
   U2430 : OAI22_X1 port map( A1 => n20362, A2 => n19996, B1 => n20014, B2 => 
                           n1935, ZN => n8369);
   U2431 : OAI22_X1 port map( A1 => n20365, A2 => n19998, B1 => n20014, B2 => 
                           n1934, ZN => n8370);
   U2432 : NAND4_X1 port map( A1 => n11566, A2 => n11567, A3 => n11568, A4 => 
                           n11569, ZN => n2225);
   U2433 : XNOR2_X1 port map( A => N113, B => N148, ZN => n11568);
   U2434 : XNOR2_X1 port map( A => N115, B => N150, ZN => n11567);
   U2435 : INV_X1 port map( A => N149, ZN => n1947);
   U2436 : NAND2_X1 port map( A1 => n11684, A2 => n11673, ZN => n3150);
   U2437 : NAND2_X1 port map( A1 => n11673, A2 => n11670, ZN => n3155);
   U2438 : AND3_X1 port map( A1 => n11672, A2 => n1939, A3 => n11688, ZN => 
                           n11676);
   U2439 : XNOR2_X1 port map( A => n11740, B => n11728, ZN => n11743);
   U2440 : AND3_X1 port map( A1 => n11680, A2 => n11676, A3 => n11675, ZN => 
                           n3153);
   U2441 : INV_X1 port map( A => n2092, ZN => n2219);
   U2442 : INV_X1 port map( A => N150, ZN => n2207);
   U2443 : INV_X1 port map( A => N80, ZN => n11565);
   U2444 : INV_X1 port map( A => n11752, ZN => U3_U2_Z_0);
   U2445 : INV_X1 port map( A => n11751, ZN => U3_U6_Z_0);
   U2446 : INV_X1 port map( A => n11622, ZN => U3_U4_Z_0);
   U2447 : AND2_X1 port map( A1 => n11691, A2 => n11679, ZN => n3163);
   U2448 : AND2_X1 port map( A1 => n11677, A2 => n11691, ZN => n3165);
   U2449 : AND2_X1 port map( A1 => n11673, A2 => n11679, ZN => n3154);
   U2450 : AND2_X1 port map( A1 => n11705, A2 => n11679, ZN => n3180);
   U2451 : INV_X1 port map( A => n11717, ZN => n3190);
   U2452 : AOI22_X1 port map( A1 => n11706, A2 => n11691, B1 => n2216, B2 => 
                           n11711, ZN => n11717);
   U2453 : AND2_X1 port map( A1 => n11705, A2 => n11706, ZN => n3184);
   U2454 : INV_X1 port map( A => n1871, ZN => n1943);
   U2455 : INV_X1 port map( A => N79, ZN => n11660);
   U2456 : INV_X1 port map( A => n11739, ZN => n11736);
   U2457 : INV_X1 port map( A => n11729, ZN => n11723);
   U2458 : OR3_X1 port map( A1 => n11671, A2 => n1939, A3 => n11672, ZN => 
                           n11699);
   U2459 : AND4_X1 port map( A1 => n2225, A2 => n11556, A3 => n2222, A4 => 
                           n2231, ZN => n2252);
   U2460 : AND4_X1 port map( A1 => n2222, A2 => n2225, A3 => n2228, A4 => n2231
                           , ZN => n2087);
   U2461 : INV_X1 port map( A => N114, ZN => n11621);
   U2462 : INV_X1 port map( A => N115, ZN => n11616);
   U2463 : INV_X1 port map( A => n11731, ZN => n11735);
   U2464 : OAI221_X1 port map( B1 => n1869, B2 => n2014, C1 => n1868, C2 => 
                           n2015, A => n20354, ZN => n2377);
   U2465 : OAI221_X1 port map( B1 => n1869, B2 => n2085, C1 => n1868, C2 => 
                           n2086, A => n20354, ZN => n2766);
   U2466 : INV_X1 port map( A => n18902, ZN => n18915);
   U2467 : INV_X1 port map( A => n18902, ZN => n18917);
   U2468 : INV_X1 port map( A => n18902, ZN => n18916);
   U2469 : BUF_X1 port map( A => n2770, Z => n19481);
   U2470 : BUF_X1 port map( A => n2770, Z => n19482);
   U2471 : BUF_X1 port map( A => n2771, Z => n19475);
   U2472 : BUF_X1 port map( A => n2771, Z => n19476);
   U2473 : BUF_X1 port map( A => n3033, Z => n19265);
   U2474 : BUF_X1 port map( A => n3033, Z => n19264);
   U2475 : BUF_X1 port map( A => n3033, Z => n19263);
   U2476 : BUF_X1 port map( A => n3033, Z => n19262);
   U2477 : INV_X1 port map( A => N113, ZN => n11613);
   U2478 : BUF_X1 port map( A => n2770, Z => n19479);
   U2479 : BUF_X1 port map( A => n2770, Z => n19480);
   U2480 : BUF_X1 port map( A => n2770, Z => n19478);
   U2481 : BUF_X1 port map( A => n2771, Z => n19473);
   U2482 : BUF_X1 port map( A => n2771, Z => n19474);
   U2483 : BUF_X1 port map( A => n2771, Z => n19472);
   U2484 : BUF_X1 port map( A => n1701, Z => n20352);
   U2485 : INV_X1 port map( A => N78, ZN => n11655);
   U2486 : BUF_X1 port map( A => n1660, Z => n20463);
   U2487 : BUF_X1 port map( A => n1659, Z => n20466);
   U2488 : BUF_X1 port map( A => n1658, Z => n20469);
   U2489 : BUF_X1 port map( A => n1657, Z => n20472);
   U2490 : BUF_X1 port map( A => n1656, Z => n20475);
   U2491 : BUF_X1 port map( A => n1655, Z => n20478);
   U2492 : BUF_X1 port map( A => n1654, Z => n20481);
   U2493 : BUF_X1 port map( A => n1653, Z => n20484);
   U2494 : BUF_X1 port map( A => n1652, Z => n20487);
   U2495 : BUF_X1 port map( A => n1651, Z => n20490);
   U2496 : BUF_X1 port map( A => n1650, Z => n20493);
   U2497 : BUF_X1 port map( A => n1649, Z => n20496);
   U2498 : BUF_X1 port map( A => n1648, Z => n20499);
   U2499 : BUF_X1 port map( A => n1647, Z => n20502);
   U2500 : BUF_X1 port map( A => n1646, Z => n20505);
   U2501 : BUF_X1 port map( A => n1645, Z => n20508);
   U2502 : BUF_X1 port map( A => n1644, Z => n20511);
   U2503 : BUF_X1 port map( A => n1643, Z => n20514);
   U2504 : BUF_X1 port map( A => n1642, Z => n20517);
   U2505 : BUF_X1 port map( A => n1641, Z => n20520);
   U2506 : BUF_X1 port map( A => n1640, Z => n20523);
   U2507 : BUF_X1 port map( A => n1639, Z => n20526);
   U2508 : BUF_X1 port map( A => n1638, Z => n20529);
   U2509 : BUF_X1 port map( A => n1637, Z => n20532);
   U2510 : BUF_X1 port map( A => n1636, Z => n20535);
   U2511 : BUF_X1 port map( A => n1635, Z => n20538);
   U2512 : BUF_X1 port map( A => n1634, Z => n20541);
   U2513 : BUF_X1 port map( A => n1631, Z => n20572);
   U2514 : BUF_X1 port map( A => n1692, Z => n20367);
   U2515 : BUF_X1 port map( A => n1691, Z => n20370);
   U2516 : BUF_X1 port map( A => n1690, Z => n20373);
   U2517 : BUF_X1 port map( A => n1689, Z => n20376);
   U2518 : BUF_X1 port map( A => n1688, Z => n20379);
   U2519 : BUF_X1 port map( A => n1687, Z => n20382);
   U2520 : BUF_X1 port map( A => n1686, Z => n20385);
   U2521 : BUF_X1 port map( A => n1685, Z => n20388);
   U2522 : BUF_X1 port map( A => n1684, Z => n20391);
   U2523 : BUF_X1 port map( A => n1683, Z => n20394);
   U2524 : BUF_X1 port map( A => n1682, Z => n20397);
   U2525 : BUF_X1 port map( A => n1681, Z => n20400);
   U2526 : BUF_X1 port map( A => n1680, Z => n20403);
   U2527 : BUF_X1 port map( A => n1679, Z => n20406);
   U2528 : BUF_X1 port map( A => n1678, Z => n20409);
   U2529 : BUF_X1 port map( A => n1677, Z => n20412);
   U2530 : BUF_X1 port map( A => n1676, Z => n20415);
   U2531 : BUF_X1 port map( A => n1675, Z => n20418);
   U2532 : BUF_X1 port map( A => n1674, Z => n20421);
   U2533 : BUF_X1 port map( A => n1673, Z => n20424);
   U2534 : BUF_X1 port map( A => n1672, Z => n20427);
   U2535 : BUF_X1 port map( A => n1671, Z => n20430);
   U2536 : BUF_X1 port map( A => n1670, Z => n20433);
   U2537 : BUF_X1 port map( A => n1669, Z => n20436);
   U2538 : BUF_X1 port map( A => n1668, Z => n20439);
   U2539 : BUF_X1 port map( A => n1667, Z => n20442);
   U2540 : BUF_X1 port map( A => n1666, Z => n20445);
   U2541 : BUF_X1 port map( A => n1665, Z => n20448);
   U2542 : BUF_X1 port map( A => n1664, Z => n20451);
   U2543 : BUF_X1 port map( A => n1663, Z => n20454);
   U2544 : BUF_X1 port map( A => n1662, Z => n20457);
   U2545 : BUF_X1 port map( A => n1661, Z => n20460);
   U2546 : BUF_X1 port map( A => n1695, Z => n20358);
   U2547 : BUF_X1 port map( A => n1694, Z => n20361);
   U2548 : BUF_X1 port map( A => n1693, Z => n20364);
   U2549 : BUF_X1 port map( A => n1660, Z => n20464);
   U2550 : BUF_X1 port map( A => n1659, Z => n20467);
   U2551 : BUF_X1 port map( A => n1658, Z => n20470);
   U2552 : BUF_X1 port map( A => n1657, Z => n20473);
   U2553 : BUF_X1 port map( A => n1656, Z => n20476);
   U2554 : BUF_X1 port map( A => n1655, Z => n20479);
   U2555 : BUF_X1 port map( A => n1654, Z => n20482);
   U2556 : BUF_X1 port map( A => n1653, Z => n20485);
   U2557 : BUF_X1 port map( A => n1652, Z => n20488);
   U2558 : BUF_X1 port map( A => n1651, Z => n20491);
   U2559 : BUF_X1 port map( A => n1650, Z => n20494);
   U2560 : BUF_X1 port map( A => n1649, Z => n20497);
   U2561 : BUF_X1 port map( A => n1648, Z => n20500);
   U2562 : BUF_X1 port map( A => n1647, Z => n20503);
   U2563 : BUF_X1 port map( A => n1646, Z => n20506);
   U2564 : BUF_X1 port map( A => n1645, Z => n20509);
   U2565 : BUF_X1 port map( A => n1644, Z => n20512);
   U2566 : BUF_X1 port map( A => n1643, Z => n20515);
   U2567 : BUF_X1 port map( A => n1642, Z => n20518);
   U2568 : BUF_X1 port map( A => n1641, Z => n20521);
   U2569 : BUF_X1 port map( A => n1640, Z => n20524);
   U2570 : BUF_X1 port map( A => n1639, Z => n20527);
   U2571 : BUF_X1 port map( A => n1638, Z => n20530);
   U2572 : BUF_X1 port map( A => n1637, Z => n20533);
   U2573 : BUF_X1 port map( A => n1636, Z => n20536);
   U2574 : BUF_X1 port map( A => n1635, Z => n20539);
   U2575 : BUF_X1 port map( A => n1634, Z => n20542);
   U2576 : BUF_X1 port map( A => n1631, Z => n20573);
   U2577 : BUF_X1 port map( A => n1692, Z => n20368);
   U2578 : BUF_X1 port map( A => n1691, Z => n20371);
   U2579 : BUF_X1 port map( A => n1690, Z => n20374);
   U2580 : BUF_X1 port map( A => n1689, Z => n20377);
   U2581 : BUF_X1 port map( A => n1688, Z => n20380);
   U2582 : BUF_X1 port map( A => n1687, Z => n20383);
   U2583 : BUF_X1 port map( A => n1686, Z => n20386);
   U2584 : BUF_X1 port map( A => n1685, Z => n20389);
   U2585 : BUF_X1 port map( A => n1684, Z => n20392);
   U2586 : BUF_X1 port map( A => n1683, Z => n20395);
   U2587 : BUF_X1 port map( A => n1682, Z => n20398);
   U2588 : BUF_X1 port map( A => n1681, Z => n20401);
   U2589 : BUF_X1 port map( A => n1680, Z => n20404);
   U2590 : BUF_X1 port map( A => n1679, Z => n20407);
   U2591 : BUF_X1 port map( A => n1678, Z => n20410);
   U2592 : BUF_X1 port map( A => n1677, Z => n20413);
   U2593 : BUF_X1 port map( A => n1676, Z => n20416);
   U2594 : BUF_X1 port map( A => n1675, Z => n20419);
   U2595 : BUF_X1 port map( A => n1674, Z => n20422);
   U2596 : BUF_X1 port map( A => n1673, Z => n20425);
   U2597 : BUF_X1 port map( A => n1672, Z => n20428);
   U2598 : BUF_X1 port map( A => n1671, Z => n20431);
   U2599 : BUF_X1 port map( A => n1670, Z => n20434);
   U2600 : BUF_X1 port map( A => n1669, Z => n20437);
   U2601 : BUF_X1 port map( A => n1668, Z => n20440);
   U2602 : BUF_X1 port map( A => n1667, Z => n20443);
   U2603 : BUF_X1 port map( A => n1666, Z => n20446);
   U2604 : BUF_X1 port map( A => n1665, Z => n20449);
   U2605 : BUF_X1 port map( A => n1664, Z => n20452);
   U2606 : BUF_X1 port map( A => n1663, Z => n20455);
   U2607 : BUF_X1 port map( A => n1662, Z => n20458);
   U2608 : BUF_X1 port map( A => n1661, Z => n20461);
   U2609 : BUF_X1 port map( A => n1696, Z => n20355);
   U2610 : BUF_X1 port map( A => n1696, Z => n20356);
   U2611 : BUF_X1 port map( A => n1695, Z => n20359);
   U2612 : BUF_X1 port map( A => n1694, Z => n20362);
   U2613 : BUF_X1 port map( A => n1693, Z => n20365);
   U2614 : BUF_X1 port map( A => n3033, Z => n19261);
   U2615 : BUF_X1 port map( A => n1660, Z => n20465);
   U2616 : BUF_X1 port map( A => n1659, Z => n20468);
   U2617 : BUF_X1 port map( A => n1658, Z => n20471);
   U2618 : BUF_X1 port map( A => n1657, Z => n20474);
   U2619 : BUF_X1 port map( A => n1656, Z => n20477);
   U2620 : BUF_X1 port map( A => n1655, Z => n20480);
   U2621 : BUF_X1 port map( A => n1654, Z => n20483);
   U2622 : BUF_X1 port map( A => n1653, Z => n20486);
   U2623 : BUF_X1 port map( A => n1652, Z => n20489);
   U2624 : BUF_X1 port map( A => n1651, Z => n20492);
   U2625 : BUF_X1 port map( A => n1650, Z => n20495);
   U2626 : BUF_X1 port map( A => n1649, Z => n20498);
   U2627 : BUF_X1 port map( A => n1648, Z => n20501);
   U2628 : BUF_X1 port map( A => n1647, Z => n20504);
   U2629 : BUF_X1 port map( A => n1646, Z => n20507);
   U2630 : BUF_X1 port map( A => n1645, Z => n20510);
   U2631 : BUF_X1 port map( A => n1644, Z => n20513);
   U2632 : BUF_X1 port map( A => n1643, Z => n20516);
   U2633 : BUF_X1 port map( A => n1642, Z => n20519);
   U2634 : BUF_X1 port map( A => n1641, Z => n20522);
   U2635 : BUF_X1 port map( A => n1640, Z => n20525);
   U2636 : BUF_X1 port map( A => n1639, Z => n20528);
   U2637 : BUF_X1 port map( A => n1638, Z => n20531);
   U2638 : BUF_X1 port map( A => n1637, Z => n20534);
   U2639 : BUF_X1 port map( A => n1636, Z => n20537);
   U2640 : BUF_X1 port map( A => n1635, Z => n20540);
   U2641 : BUF_X1 port map( A => n1634, Z => n20543);
   U2642 : BUF_X1 port map( A => n1631, Z => n20574);
   U2643 : BUF_X1 port map( A => n1692, Z => n20369);
   U2644 : BUF_X1 port map( A => n1691, Z => n20372);
   U2645 : BUF_X1 port map( A => n1690, Z => n20375);
   U2646 : BUF_X1 port map( A => n1689, Z => n20378);
   U2647 : BUF_X1 port map( A => n1688, Z => n20381);
   U2648 : BUF_X1 port map( A => n1687, Z => n20384);
   U2649 : BUF_X1 port map( A => n1686, Z => n20387);
   U2650 : BUF_X1 port map( A => n1685, Z => n20390);
   U2651 : BUF_X1 port map( A => n1684, Z => n20393);
   U2652 : BUF_X1 port map( A => n1683, Z => n20396);
   U2653 : BUF_X1 port map( A => n1682, Z => n20399);
   U2654 : BUF_X1 port map( A => n1681, Z => n20402);
   U2655 : BUF_X1 port map( A => n1680, Z => n20405);
   U2656 : BUF_X1 port map( A => n1679, Z => n20408);
   U2657 : BUF_X1 port map( A => n1678, Z => n20411);
   U2658 : BUF_X1 port map( A => n1677, Z => n20414);
   U2659 : BUF_X1 port map( A => n1676, Z => n20417);
   U2660 : BUF_X1 port map( A => n1675, Z => n20420);
   U2661 : BUF_X1 port map( A => n1674, Z => n20423);
   U2662 : BUF_X1 port map( A => n1673, Z => n20426);
   U2663 : BUF_X1 port map( A => n1672, Z => n20429);
   U2664 : BUF_X1 port map( A => n1671, Z => n20432);
   U2665 : BUF_X1 port map( A => n1670, Z => n20435);
   U2666 : BUF_X1 port map( A => n1669, Z => n20438);
   U2667 : BUF_X1 port map( A => n1668, Z => n20441);
   U2668 : BUF_X1 port map( A => n1667, Z => n20444);
   U2669 : BUF_X1 port map( A => n1666, Z => n20447);
   U2670 : BUF_X1 port map( A => n1665, Z => n20450);
   U2671 : BUF_X1 port map( A => n1664, Z => n20453);
   U2672 : BUF_X1 port map( A => n1663, Z => n20456);
   U2673 : BUF_X1 port map( A => n1662, Z => n20459);
   U2674 : BUF_X1 port map( A => n1661, Z => n20462);
   U2675 : BUF_X1 port map( A => n1696, Z => n20357);
   U2676 : BUF_X1 port map( A => n1695, Z => n20360);
   U2677 : BUF_X1 port map( A => n1694, Z => n20363);
   U2678 : BUF_X1 port map( A => n1693, Z => n20366);
   U2679 : BUF_X1 port map( A => n1701, Z => n20353);
   U2680 : BUF_X1 port map( A => n1701, Z => n20354);
   U2681 : INV_X1 port map( A => n11680, ZN => n11674);
   U2682 : XNOR2_X1 port map( A => count3(2), B => n11731, ZN => n11755);
   U2683 : OAI211_X1 port map( C1 => n11739, C2 => n11740, A => n11741, B => 
                           n11726, ZN => n11672);
   U2684 : OAI21_X1 port map( B1 => n11742, B2 => n11736, A => count3(3), ZN =>
                           n11741);
   U2685 : INV_X1 port map( A => n11740, ZN => n11742);
   U2686 : XNOR2_X1 port map( A => n11724, B => count3(3), ZN => n11722);
   U2687 : NOR3_X1 port map( A1 => n11688, A2 => count3(0), A3 => n11672, ZN =>
                           n11691);
   U2688 : AOI21_X1 port map( B1 => add_rd2(3), B2 => n11757, A => add_rd2(4), 
                           ZN => n11622);
   U2689 : OR3_X1 port map( A1 => add_rd2(2), A2 => add_rd2(1), A3 => 
                           add_rd2(0), ZN => n11757);
   U2690 : OAI222_X1 port map( A1 => n3502, A2 => n19134, B1 => n2763, B2 => 
                           n19128, C1 => n3434, C2 => n19122, ZN => n11647);
   U2691 : OAI222_X1 port map( A1 => n3502, A2 => n19333, B1 => n2763, B2 => 
                           n19327, C1 => n3434, C2 => n19321, ZN => n11607);
   U2692 : OAI222_X1 port map( A1 => n3501, A2 => n19134, B1 => n2762, B2 => 
                           n19128, C1 => n3433, C2 => n19122, ZN => n11528);
   U2693 : OAI222_X1 port map( A1 => n3501, A2 => n19333, B1 => n2762, B2 => 
                           n19327, C1 => n3433, C2 => n19321, ZN => n11508);
   U2694 : OAI222_X1 port map( A1 => n3500, A2 => n19134, B1 => n2761, B2 => 
                           n19128, C1 => n3432, C2 => n19122, ZN => n11461);
   U2695 : OAI222_X1 port map( A1 => n3500, A2 => n19333, B1 => n2761, B2 => 
                           n19327, C1 => n3432, C2 => n19321, ZN => n11441);
   U2696 : OAI222_X1 port map( A1 => n3499, A2 => n19134, B1 => n2760, B2 => 
                           n19128, C1 => n3431, C2 => n19122, ZN => n11394);
   U2697 : OAI222_X1 port map( A1 => n3499, A2 => n19333, B1 => n2760, B2 => 
                           n19327, C1 => n3431, C2 => n19321, ZN => n11373);
   U2698 : OAI222_X1 port map( A1 => n3498, A2 => n19134, B1 => n2759, B2 => 
                           n19128, C1 => n3430, C2 => n19122, ZN => n11326);
   U2699 : OAI222_X1 port map( A1 => n3498, A2 => n19333, B1 => n2759, B2 => 
                           n19327, C1 => n3430, C2 => n19321, ZN => n11306);
   U2700 : OAI222_X1 port map( A1 => n3497, A2 => n19134, B1 => n2758, B2 => 
                           n19128, C1 => n3429, C2 => n19122, ZN => n11259);
   U2701 : OAI222_X1 port map( A1 => n3497, A2 => n19333, B1 => n2758, B2 => 
                           n19327, C1 => n3429, C2 => n19321, ZN => n11239);
   U2702 : OAI222_X1 port map( A1 => n3496, A2 => n19134, B1 => n2757, B2 => 
                           n19128, C1 => n3428, C2 => n19122, ZN => n11192);
   U2703 : OAI222_X1 port map( A1 => n3496, A2 => n19333, B1 => n2757, B2 => 
                           n19327, C1 => n3428, C2 => n19321, ZN => n11171);
   U2704 : OAI222_X1 port map( A1 => n3495, A2 => n19134, B1 => n2756, B2 => 
                           n19128, C1 => n3427, C2 => n19122, ZN => n11125);
   U2705 : OAI222_X1 port map( A1 => n3495, A2 => n19333, B1 => n2756, B2 => 
                           n19327, C1 => n3427, C2 => n19321, ZN => n11104);
   U2706 : OAI222_X1 port map( A1 => n3494, A2 => n19134, B1 => n2755, B2 => 
                           n19128, C1 => n3426, C2 => n19122, ZN => n11057);
   U2707 : OAI222_X1 port map( A1 => n3494, A2 => n19333, B1 => n2755, B2 => 
                           n19327, C1 => n3426, C2 => n19321, ZN => n11037);
   U2708 : OAI222_X1 port map( A1 => n3493, A2 => n19134, B1 => n2754, B2 => 
                           n19128, C1 => n3425, C2 => n19122, ZN => n10990);
   U2709 : OAI222_X1 port map( A1 => n3493, A2 => n19333, B1 => n2754, B2 => 
                           n19327, C1 => n3425, C2 => n19321, ZN => n10970);
   U2710 : OAI222_X1 port map( A1 => n3492, A2 => n19134, B1 => n2753, B2 => 
                           n19128, C1 => n3424, C2 => n19122, ZN => n10923);
   U2711 : OAI222_X1 port map( A1 => n3492, A2 => n19333, B1 => n2753, B2 => 
                           n19327, C1 => n3424, C2 => n19321, ZN => n10902);
   U2712 : OAI222_X1 port map( A1 => n3491, A2 => n19134, B1 => n2752, B2 => 
                           n19128, C1 => n3423, C2 => n19122, ZN => n10856);
   U2713 : OAI222_X1 port map( A1 => n3491, A2 => n19333, B1 => n2752, B2 => 
                           n19327, C1 => n3423, C2 => n19321, ZN => n10835);
   U2714 : OAI222_X1 port map( A1 => n3490, A2 => n19135, B1 => n2751, B2 => 
                           n19129, C1 => n3422, C2 => n19123, ZN => n10788);
   U2715 : OAI222_X1 port map( A1 => n3490, A2 => n19334, B1 => n2751, B2 => 
                           n19328, C1 => n3422, C2 => n19322, ZN => n10768);
   U2716 : OAI222_X1 port map( A1 => n3489, A2 => n19135, B1 => n2750, B2 => 
                           n19129, C1 => n3421, C2 => n19123, ZN => n10721);
   U2717 : OAI222_X1 port map( A1 => n3489, A2 => n19334, B1 => n2750, B2 => 
                           n19328, C1 => n3421, C2 => n19322, ZN => n10701);
   U2718 : OAI222_X1 port map( A1 => n3488, A2 => n19135, B1 => n2749, B2 => 
                           n19129, C1 => n3420, C2 => n19123, ZN => n10654);
   U2719 : OAI222_X1 port map( A1 => n3488, A2 => n19334, B1 => n2749, B2 => 
                           n19328, C1 => n3420, C2 => n19322, ZN => n10633);
   U2720 : OAI222_X1 port map( A1 => n3487, A2 => n19135, B1 => n2748, B2 => 
                           n19129, C1 => n3419, C2 => n19123, ZN => n10586);
   U2721 : OAI222_X1 port map( A1 => n3487, A2 => n19334, B1 => n2748, B2 => 
                           n19328, C1 => n3419, C2 => n19322, ZN => n10566);
   U2722 : OAI222_X1 port map( A1 => n3486, A2 => n19135, B1 => n2747, B2 => 
                           n19129, C1 => n3418, C2 => n19123, ZN => n10519);
   U2723 : OAI222_X1 port map( A1 => n3486, A2 => n19334, B1 => n2747, B2 => 
                           n19328, C1 => n3418, C2 => n19322, ZN => n10499);
   U2724 : OAI222_X1 port map( A1 => n3485, A2 => n19135, B1 => n2746, B2 => 
                           n19129, C1 => n3417, C2 => n19123, ZN => n10452);
   U2725 : OAI222_X1 port map( A1 => n3485, A2 => n19334, B1 => n2746, B2 => 
                           n19328, C1 => n3417, C2 => n19322, ZN => n10432);
   U2726 : OAI222_X1 port map( A1 => n3484, A2 => n19135, B1 => n2745, B2 => 
                           n19129, C1 => n3416, C2 => n19123, ZN => n10385);
   U2727 : OAI222_X1 port map( A1 => n3484, A2 => n19334, B1 => n2745, B2 => 
                           n19328, C1 => n3416, C2 => n19322, ZN => n10364);
   U2728 : OAI222_X1 port map( A1 => n3483, A2 => n19135, B1 => n2744, B2 => 
                           n19129, C1 => n3415, C2 => n19123, ZN => n10317);
   U2729 : OAI222_X1 port map( A1 => n3483, A2 => n19334, B1 => n2744, B2 => 
                           n19328, C1 => n3415, C2 => n19322, ZN => n10297);
   U2730 : OAI222_X1 port map( A1 => n3482, A2 => n19135, B1 => n2743, B2 => 
                           n19129, C1 => n3414, C2 => n19123, ZN => n10250);
   U2731 : OAI222_X1 port map( A1 => n3482, A2 => n19334, B1 => n2743, B2 => 
                           n19328, C1 => n3414, C2 => n19322, ZN => n10230);
   U2732 : OAI222_X1 port map( A1 => n3481, A2 => n19135, B1 => n2742, B2 => 
                           n19129, C1 => n3413, C2 => n19123, ZN => n10183);
   U2733 : OAI222_X1 port map( A1 => n3481, A2 => n19334, B1 => n2742, B2 => 
                           n19328, C1 => n3413, C2 => n19322, ZN => n10162);
   U2734 : OAI222_X1 port map( A1 => n3480, A2 => n19135, B1 => n2741, B2 => 
                           n19129, C1 => n3412, C2 => n19123, ZN => n10116);
   U2735 : OAI222_X1 port map( A1 => n3480, A2 => n19334, B1 => n2741, B2 => 
                           n19328, C1 => n3412, C2 => n19322, ZN => n10095);
   U2736 : OAI222_X1 port map( A1 => n3479, A2 => n19135, B1 => n2740, B2 => 
                           n19129, C1 => n3411, C2 => n19123, ZN => n10048);
   U2737 : OAI222_X1 port map( A1 => n3479, A2 => n19334, B1 => n2740, B2 => 
                           n19328, C1 => n3411, C2 => n19322, ZN => n10028);
   U2738 : OAI222_X1 port map( A1 => n3478, A2 => n19136, B1 => n2739, B2 => 
                           n19130, C1 => n3410, C2 => n19124, ZN => n9981);
   U2739 : OAI222_X1 port map( A1 => n3478, A2 => n19335, B1 => n2739, B2 => 
                           n19329, C1 => n3410, C2 => n19323, ZN => n9961);
   U2740 : OAI222_X1 port map( A1 => n3477, A2 => n19136, B1 => n2738, B2 => 
                           n19130, C1 => n3409, C2 => n19124, ZN => n9914);
   U2741 : OAI222_X1 port map( A1 => n3477, A2 => n19335, B1 => n2738, B2 => 
                           n19329, C1 => n3409, C2 => n19323, ZN => n9893);
   U2742 : OAI222_X1 port map( A1 => n3476, A2 => n19136, B1 => n2737, B2 => 
                           n19130, C1 => n3408, C2 => n19124, ZN => n9846);
   U2743 : OAI222_X1 port map( A1 => n3476, A2 => n19335, B1 => n2737, B2 => 
                           n19329, C1 => n3408, C2 => n19323, ZN => n9826);
   U2744 : OAI222_X1 port map( A1 => n3475, A2 => n19136, B1 => n2736, B2 => 
                           n19130, C1 => n3407, C2 => n19124, ZN => n9779);
   U2745 : OAI222_X1 port map( A1 => n3475, A2 => n19335, B1 => n2736, B2 => 
                           n19329, C1 => n3407, C2 => n19323, ZN => n9759);
   U2746 : OAI222_X1 port map( A1 => n3474, A2 => n19136, B1 => n2735, B2 => 
                           n19130, C1 => n3406, C2 => n19124, ZN => n9712);
   U2747 : OAI222_X1 port map( A1 => n3474, A2 => n19335, B1 => n2735, B2 => 
                           n19329, C1 => n3406, C2 => n19323, ZN => n9692);
   U2748 : OAI222_X1 port map( A1 => n3473, A2 => n19136, B1 => n2734, B2 => 
                           n19130, C1 => n3405, C2 => n19124, ZN => n9645);
   U2749 : OAI222_X1 port map( A1 => n3473, A2 => n19335, B1 => n2734, B2 => 
                           n19329, C1 => n3405, C2 => n19323, ZN => n9624);
   U2750 : OAI222_X1 port map( A1 => n3472, A2 => n19136, B1 => n2733, B2 => 
                           n19130, C1 => n3404, C2 => n19124, ZN => n9577);
   U2751 : OAI222_X1 port map( A1 => n3472, A2 => n19335, B1 => n2733, B2 => 
                           n19329, C1 => n3404, C2 => n19323, ZN => n9557);
   U2752 : OAI222_X1 port map( A1 => n3471, A2 => n19136, B1 => n2732, B2 => 
                           n19130, C1 => n3403, C2 => n19124, ZN => n9510);
   U2753 : OAI222_X1 port map( A1 => n3471, A2 => n19335, B1 => n2732, B2 => 
                           n19329, C1 => n3403, C2 => n19323, ZN => n9490);
   U2754 : OAI222_X1 port map( A1 => n3470, A2 => n19136, B1 => n2731, B2 => 
                           n19130, C1 => n3402, C2 => n19124, ZN => n9443);
   U2755 : OAI222_X1 port map( A1 => n3470, A2 => n19335, B1 => n2731, B2 => 
                           n19329, C1 => n3402, C2 => n19323, ZN => n9422);
   U2756 : OAI222_X1 port map( A1 => n3469, A2 => n19136, B1 => n2730, B2 => 
                           n19130, C1 => n3401, C2 => n19124, ZN => n9376);
   U2757 : OAI222_X1 port map( A1 => n3469, A2 => n19335, B1 => n2730, B2 => 
                           n19329, C1 => n3401, C2 => n19323, ZN => n9355);
   U2758 : OAI222_X1 port map( A1 => n3468, A2 => n19136, B1 => n2729, B2 => 
                           n19130, C1 => n3400, C2 => n19124, ZN => n9308);
   U2759 : OAI222_X1 port map( A1 => n3468, A2 => n19335, B1 => n2729, B2 => 
                           n19329, C1 => n3400, C2 => n19323, ZN => n9288);
   U2760 : OAI222_X1 port map( A1 => n3467, A2 => n19136, B1 => n2728, B2 => 
                           n19130, C1 => n3399, C2 => n19124, ZN => n7001);
   U2761 : OAI222_X1 port map( A1 => n3467, A2 => n19335, B1 => n2728, B2 => 
                           n19329, C1 => n3399, C2 => n19323, ZN => n6981);
   U2762 : OAI222_X1 port map( A1 => n3466, A2 => n19137, B1 => n2727, B2 => 
                           n19131, C1 => n3398, C2 => n19125, ZN => n6934);
   U2763 : OAI222_X1 port map( A1 => n3466, A2 => n19336, B1 => n2727, B2 => 
                           n19330, C1 => n3398, C2 => n19324, ZN => n6914);
   U2764 : OAI222_X1 port map( A1 => n3465, A2 => n19137, B1 => n2726, B2 => 
                           n19131, C1 => n3397, C2 => n19125, ZN => n6868);
   U2765 : OAI222_X1 port map( A1 => n3465, A2 => n19336, B1 => n2726, B2 => 
                           n19330, C1 => n3397, C2 => n19324, ZN => n6847);
   U2766 : OAI222_X1 port map( A1 => n3464, A2 => n19137, B1 => n2725, B2 => 
                           n19131, C1 => n3396, C2 => n19125, ZN => n6800);
   U2767 : OAI222_X1 port map( A1 => n3464, A2 => n19336, B1 => n2725, B2 => 
                           n19330, C1 => n3396, C2 => n19324, ZN => n6780);
   U2768 : OAI222_X1 port map( A1 => n3463, A2 => n19137, B1 => n2724, B2 => 
                           n19131, C1 => n3395, C2 => n19125, ZN => n6733);
   U2769 : OAI222_X1 port map( A1 => n3463, A2 => n19336, B1 => n2724, B2 => 
                           n19330, C1 => n3395, C2 => n19324, ZN => n6713);
   U2770 : OAI222_X1 port map( A1 => n3462, A2 => n19137, B1 => n2723, B2 => 
                           n19131, C1 => n3394, C2 => n19125, ZN => n6666);
   U2771 : OAI222_X1 port map( A1 => n3462, A2 => n19336, B1 => n2723, B2 => 
                           n19330, C1 => n3394, C2 => n19324, ZN => n6646);
   U2772 : OAI222_X1 port map( A1 => n3461, A2 => n19137, B1 => n2722, B2 => 
                           n19131, C1 => n3393, C2 => n19125, ZN => n6599);
   U2773 : OAI222_X1 port map( A1 => n3461, A2 => n19336, B1 => n2722, B2 => 
                           n19330, C1 => n3393, C2 => n19324, ZN => n6579);
   U2774 : OAI222_X1 port map( A1 => n3460, A2 => n19137, B1 => n2721, B2 => 
                           n19131, C1 => n3392, C2 => n19125, ZN => n6533);
   U2775 : OAI222_X1 port map( A1 => n3460, A2 => n19336, B1 => n2721, B2 => 
                           n19330, C1 => n3392, C2 => n19324, ZN => n6513);
   U2776 : OAI222_X1 port map( A1 => n3459, A2 => n19137, B1 => n2720, B2 => 
                           n19131, C1 => n3391, C2 => n19125, ZN => n6467);
   U2777 : OAI222_X1 port map( A1 => n3459, A2 => n19336, B1 => n2720, B2 => 
                           n19330, C1 => n3391, C2 => n19324, ZN => n6447);
   U2778 : OAI222_X1 port map( A1 => n3458, A2 => n19137, B1 => n2463, B2 => 
                           n19131, C1 => n3390, C2 => n19125, ZN => n6401);
   U2779 : OAI222_X1 port map( A1 => n3458, A2 => n19336, B1 => n2463, B2 => 
                           n19330, C1 => n3390, C2 => n19324, ZN => n6381);
   U2780 : OAI222_X1 port map( A1 => n3457, A2 => n19137, B1 => n2462, B2 => 
                           n19131, C1 => n3389, C2 => n19125, ZN => n6335);
   U2781 : OAI222_X1 port map( A1 => n3457, A2 => n19336, B1 => n2462, B2 => 
                           n19330, C1 => n3389, C2 => n19324, ZN => n6315);
   U2782 : OAI222_X1 port map( A1 => n3456, A2 => n19137, B1 => n2461, B2 => 
                           n19131, C1 => n3388, C2 => n19125, ZN => n6269);
   U2783 : OAI222_X1 port map( A1 => n3456, A2 => n19336, B1 => n2461, B2 => 
                           n19330, C1 => n3388, C2 => n19324, ZN => n6249);
   U2784 : OAI222_X1 port map( A1 => n3455, A2 => n19137, B1 => n2460, B2 => 
                           n19131, C1 => n3387, C2 => n19125, ZN => n6203);
   U2785 : OAI222_X1 port map( A1 => n3455, A2 => n19336, B1 => n2460, B2 => 
                           n19330, C1 => n3387, C2 => n19324, ZN => n6183);
   U2786 : OAI222_X1 port map( A1 => n3454, A2 => n19138, B1 => n2459, B2 => 
                           n19132, C1 => n3386, C2 => n19126, ZN => n6137);
   U2787 : OAI222_X1 port map( A1 => n3454, A2 => n19337, B1 => n2459, B2 => 
                           n19331, C1 => n3386, C2 => n19325, ZN => n6117);
   U2788 : OAI222_X1 port map( A1 => n3453, A2 => n19138, B1 => n2458, B2 => 
                           n19132, C1 => n3385, C2 => n19126, ZN => n6071);
   U2789 : OAI222_X1 port map( A1 => n3453, A2 => n19337, B1 => n2458, B2 => 
                           n19331, C1 => n3385, C2 => n19325, ZN => n6051);
   U2790 : OAI222_X1 port map( A1 => n3452, A2 => n19138, B1 => n2457, B2 => 
                           n19132, C1 => n3384, C2 => n19126, ZN => n6003);
   U2791 : OAI222_X1 port map( A1 => n3452, A2 => n19337, B1 => n2457, B2 => 
                           n19331, C1 => n3384, C2 => n19325, ZN => n5983);
   U2792 : OAI222_X1 port map( A1 => n3451, A2 => n19138, B1 => n2456, B2 => 
                           n19132, C1 => n3383, C2 => n19126, ZN => n5935);
   U2793 : OAI222_X1 port map( A1 => n3451, A2 => n19337, B1 => n2456, B2 => 
                           n19331, C1 => n3383, C2 => n19325, ZN => n5915);
   U2794 : OAI222_X1 port map( A1 => n3450, A2 => n19138, B1 => n2455, B2 => 
                           n19132, C1 => n3382, C2 => n19126, ZN => n5868);
   U2795 : OAI222_X1 port map( A1 => n3450, A2 => n19337, B1 => n2455, B2 => 
                           n19331, C1 => n3382, C2 => n19325, ZN => n5848);
   U2796 : OAI222_X1 port map( A1 => n3449, A2 => n19138, B1 => n2454, B2 => 
                           n19132, C1 => n3381, C2 => n19126, ZN => n5801);
   U2797 : OAI222_X1 port map( A1 => n3449, A2 => n19337, B1 => n2454, B2 => 
                           n19331, C1 => n3381, C2 => n19325, ZN => n5781);
   U2798 : OAI222_X1 port map( A1 => n3448, A2 => n19138, B1 => n2453, B2 => 
                           n19132, C1 => n3380, C2 => n19126, ZN => n5729);
   U2799 : OAI222_X1 port map( A1 => n3448, A2 => n19337, B1 => n2453, B2 => 
                           n19331, C1 => n3380, C2 => n19325, ZN => n5709);
   U2800 : OAI222_X1 port map( A1 => n3447, A2 => n19138, B1 => n2452, B2 => 
                           n19132, C1 => n3379, C2 => n19126, ZN => n5659);
   U2801 : OAI222_X1 port map( A1 => n3447, A2 => n19337, B1 => n2452, B2 => 
                           n19331, C1 => n3379, C2 => n19325, ZN => n5639);
   U2802 : OAI222_X1 port map( A1 => n3446, A2 => n19138, B1 => n2451, B2 => 
                           n19132, C1 => n3378, C2 => n19126, ZN => n5591);
   U2803 : OAI222_X1 port map( A1 => n3446, A2 => n19337, B1 => n2451, B2 => 
                           n19331, C1 => n3378, C2 => n19325, ZN => n5571);
   U2804 : OAI222_X1 port map( A1 => n3445, A2 => n19138, B1 => n2450, B2 => 
                           n19132, C1 => n3377, C2 => n19126, ZN => n5522);
   U2805 : OAI222_X1 port map( A1 => n3445, A2 => n19337, B1 => n2450, B2 => 
                           n19331, C1 => n3377, C2 => n19325, ZN => n5502);
   U2806 : OAI222_X1 port map( A1 => n3444, A2 => n19138, B1 => n2449, B2 => 
                           n19132, C1 => n3376, C2 => n19126, ZN => n5453);
   U2807 : OAI222_X1 port map( A1 => n3444, A2 => n19337, B1 => n2449, B2 => 
                           n19331, C1 => n3376, C2 => n19325, ZN => n5433);
   U2808 : OAI222_X1 port map( A1 => n3443, A2 => n19138, B1 => n2448, B2 => 
                           n19132, C1 => n3375, C2 => n19126, ZN => n5385);
   U2809 : OAI222_X1 port map( A1 => n3443, A2 => n19337, B1 => n2448, B2 => 
                           n19331, C1 => n3375, C2 => n19325, ZN => n5365);
   U2810 : OAI222_X1 port map( A1 => n3442, A2 => n19139, B1 => n2447, B2 => 
                           n19133, C1 => n3374, C2 => n19127, ZN => n5315);
   U2811 : OAI222_X1 port map( A1 => n3442, A2 => n19338, B1 => n2447, B2 => 
                           n19332, C1 => n3374, C2 => n19326, ZN => n5295);
   U2812 : OAI222_X1 port map( A1 => n3441, A2 => n19139, B1 => n2446, B2 => 
                           n19133, C1 => n3373, C2 => n19127, ZN => n4446);
   U2813 : OAI222_X1 port map( A1 => n3441, A2 => n19338, B1 => n2446, B2 => 
                           n19332, C1 => n3373, C2 => n19326, ZN => n4106);
   U2814 : OAI222_X1 port map( A1 => n3440, A2 => n19139, B1 => n2445, B2 => 
                           n19133, C1 => n3372, C2 => n19127, ZN => n3288);
   U2815 : OAI222_X1 port map( A1 => n3440, A2 => n19338, B1 => n2445, B2 => 
                           n19332, C1 => n3372, C2 => n19326, ZN => n3248);
   U2816 : OAI222_X1 port map( A1 => n3439, A2 => n19139, B1 => n2444, B2 => 
                           n19133, C1 => n3371, C2 => n19127, ZN => n3116);
   U2817 : OAI222_X1 port map( A1 => n3439, A2 => n19338, B1 => n2444, B2 => 
                           n19332, C1 => n3371, C2 => n19326, ZN => n2999);
   U2818 : NOR4_X1 port map( A1 => n5325, A2 => n5326, A3 => n5327, A4 => n5328
                           , ZN => n5324);
   U2819 : OAI222_X1 port map( A1 => n1733, A2 => n19073, B1 => n3776, B2 => 
                           n19067, C1 => n3710, C2 => n19061, ZN => n5328);
   U2820 : OAI221_X1 port map( B1 => n4182, B2 => n19031, C1 => n1877, C2 => 
                           n19025, A => n5330, ZN => n5326);
   U2821 : OAI221_X1 port map( B1 => n19007, B2 => n4856, C1 => n2100, C2 => 
                           n19001, A => n5331, ZN => n5325);
   U2822 : NOR4_X1 port map( A1 => n4584, A2 => n4585, A3 => n4586, A4 => n4587
                           , ZN => n4583);
   U2823 : OAI222_X1 port map( A1 => n1732, A2 => n19073, B1 => n3775, B2 => 
                           n19067, C1 => n3709, C2 => n19061, ZN => n4587);
   U2824 : OAI221_X1 port map( B1 => n4181, B2 => n19031, C1 => n1876, C2 => 
                           n19025, A => n4653, ZN => n4585);
   U2825 : OAI221_X1 port map( B1 => n19007, B2 => n3638, C1 => n2099, C2 => 
                           n19001, A => n4718, ZN => n4584);
   U2826 : NOR4_X1 port map( A1 => n3302, A2 => n3367, A3 => n3368, A4 => n3369
                           , ZN => n3301);
   U2827 : OAI222_X1 port map( A1 => n1731, A2 => n19073, B1 => n3774, B2 => 
                           n19067, C1 => n3708, C2 => n19061, ZN => n3369);
   U2828 : OAI221_X1 port map( B1 => n4180, B2 => n19031, C1 => n1875, C2 => 
                           n19025, A => n3435, ZN => n3367);
   U2829 : OAI221_X1 port map( B1 => n19007, B2 => n3208, C1 => n2098, C2 => 
                           n19001, A => n3436, ZN => n3302);
   U2830 : NOR4_X1 port map( A1 => n3143, A2 => n3144, A3 => n3145, A4 => n3146
                           , ZN => n3142);
   U2831 : OAI222_X1 port map( A1 => n1730, A2 => n19073, B1 => n3773, B2 => 
                           n19067, C1 => n3707, C2 => n19061, ZN => n3146);
   U2832 : OAI221_X1 port map( B1 => n4179, B2 => n19031, C1 => n1874, C2 => 
                           n19025, A => n3157, ZN => n3144);
   U2833 : OAI221_X1 port map( B1 => n19007, B2 => n2768, C1 => n2097, C2 => 
                           n19001, A => n3162, ZN => n3143);
   U2834 : NOR4_X1 port map( A1 => n5307, A2 => n5308, A3 => n5309, A4 => n5310
                           , ZN => n5306);
   U2835 : OAI221_X1 port map( B1 => n1877, B2 => n19272, C1 => n19261, C2 => 
                           n2325, A => n5311, ZN => n5310);
   U2836 : OAI221_X1 port map( B1 => n4861, B2 => n19248, C1 => n2381, C2 => 
                           n19242, A => n5312, ZN => n5309);
   U2837 : OAI221_X1 port map( B1 => n1803, B2 => n19200, C1 => n4182, C2 => 
                           n19194, A => n5314, ZN => n5307);
   U2838 : NOR4_X1 port map( A1 => n4989, A2 => n5054, A3 => n5055, A4 => n5056
                           , ZN => n4988);
   U2839 : OAI221_X1 port map( B1 => n1803, B2 => n19399, C1 => n4182, C2 => 
                           n19393, A => n5292, ZN => n4989);
   U2840 : OAI221_X1 port map( B1 => n1877, B2 => n19471, C1 => n19460, C2 => 
                           n2326, A => n5121, ZN => n5056);
   U2841 : OAI221_X1 port map( B1 => n4861, B2 => n19447, C1 => n2381, C2 => 
                           n19441, A => n5188, ZN => n5055);
   U2842 : NOR4_X1 port map( A1 => n4310, A2 => n4311, A3 => n4312, A4 => n4377
                           , ZN => n4245);
   U2843 : OAI221_X1 port map( B1 => n1876, B2 => n19272, C1 => n19261, C2 => 
                           n2328, A => n4378, ZN => n4377);
   U2844 : OAI221_X1 port map( B1 => n4860, B2 => n19248, C1 => n2380, C2 => 
                           n19242, A => n4379, ZN => n4312);
   U2845 : OAI221_X1 port map( B1 => n1802, B2 => n19200, C1 => n4181, C2 => 
                           n19194, A => n4445, ZN => n4310);
   U2846 : NOR4_X1 port map( A1 => n3771, A2 => n3772, A3 => n3837, A4 => n3838
                           , ZN => n3706);
   U2847 : OAI221_X1 port map( B1 => n1802, B2 => n19399, C1 => n4181, C2 => 
                           n19393, A => n4039, ZN => n3771);
   U2848 : OAI221_X1 port map( B1 => n1876, B2 => n19471, C1 => n19460, C2 => 
                           n2329, A => n3839, ZN => n3838);
   U2849 : OAI221_X1 port map( B1 => n4860, B2 => n19447, C1 => n2380, C2 => 
                           n19441, A => n3906, ZN => n3837);
   U2850 : NOR4_X1 port map( A1 => n3272, A2 => n3274, A3 => n3276, A4 => n3278
                           , ZN => n3270);
   U2851 : OAI221_X1 port map( B1 => n1875, B2 => n19272, C1 => n19261, C2 => 
                           n2331, A => n3280, ZN => n3278);
   U2852 : OAI221_X1 port map( B1 => n4859, B2 => n19248, C1 => n2379, C2 => 
                           n19242, A => n3282, ZN => n3276);
   U2853 : OAI221_X1 port map( B1 => n1801, B2 => n19200, C1 => n4180, C2 => 
                           n19194, A => n3286, ZN => n3272);
   U2854 : NOR4_X1 port map( A1 => n3218, A2 => n3220, A3 => n3222, A4 => n3224
                           , ZN => n3216);
   U2855 : OAI221_X1 port map( B1 => n1801, B2 => n19399, C1 => n4180, C2 => 
                           n19393, A => n3242, ZN => n3218);
   U2856 : OAI221_X1 port map( B1 => n1875, B2 => n19471, C1 => n19460, C2 => 
                           n2332, A => n3226, ZN => n3224);
   U2857 : OAI221_X1 port map( B1 => n4859, B2 => n19447, C1 => n2379, C2 => 
                           n19441, A => n3232, ZN => n3222);
   U2858 : NOR4_X1 port map( A1 => n3028, A2 => n3029, A3 => n3030, A4 => n3031
                           , ZN => n3027);
   U2859 : OAI221_X1 port map( B1 => n1874, B2 => n19272, C1 => n19261, C2 => 
                           n2334, A => n3034, ZN => n3031);
   U2860 : OAI221_X1 port map( B1 => n4858, B2 => n19248, C1 => n2378, C2 => 
                           n19242, A => n3103, ZN => n3030);
   U2861 : OAI221_X1 port map( B1 => n1800, B2 => n19200, C1 => n4179, C2 => 
                           n19194, A => n3113, ZN => n3028);
   U2862 : NOR4_X1 port map( A1 => n2776, A2 => n2777, A3 => n2778, A4 => n2779
                           , ZN => n2775);
   U2863 : OAI221_X1 port map( B1 => n1800, B2 => n19399, C1 => n4179, C2 => 
                           n19393, A => n2994, ZN => n2776);
   U2864 : OAI221_X1 port map( B1 => n1874, B2 => n19471, C1 => n19460, C2 => 
                           n2335, A => n2782, ZN => n2779);
   U2865 : OAI221_X1 port map( B1 => n4858, B2 => n19447, C1 => n2378, C2 => 
                           n19441, A => n2981, ZN => n2778);
   U2866 : NOR4_X1 port map( A1 => n6743, A2 => n6744, A3 => n6745, A4 => n6746
                           , ZN => n6742);
   U2867 : OAI222_X1 port map( A1 => n1757, A2 => n19071, B1 => n3797, B2 => 
                           n19065, C1 => n3731, C2 => n19059, ZN => n6746);
   U2868 : OAI221_X1 port map( B1 => n4203, B2 => n19029, C1 => n1898, C2 => 
                           n19023, A => n6748, ZN => n6744);
   U2869 : OAI221_X1 port map( B1 => n19005, B2 => n6692, C1 => n2121, C2 => 
                           n18999, A => n6750, ZN => n6743);
   U2870 : NOR4_X1 port map( A1 => n6676, A2 => n6677, A3 => n6678, A4 => n6679
                           , ZN => n6675);
   U2871 : OAI222_X1 port map( A1 => n1756, A2 => n19071, B1 => n3796, B2 => 
                           n19065, C1 => n3730, C2 => n19059, ZN => n6679);
   U2872 : OAI221_X1 port map( B1 => n4202, B2 => n19029, C1 => n1897, C2 => 
                           n19023, A => n6681, ZN => n6677);
   U2873 : OAI221_X1 port map( B1 => n19005, B2 => n6625, C1 => n2120, C2 => 
                           n18999, A => n6682, ZN => n6676);
   U2874 : NOR4_X1 port map( A1 => n6609, A2 => n6610, A3 => n6611, A4 => n6612
                           , ZN => n6608);
   U2875 : OAI222_X1 port map( A1 => n1755, A2 => n19071, B1 => n3795, B2 => 
                           n19065, C1 => n3729, C2 => n19059, ZN => n6612);
   U2876 : OAI221_X1 port map( B1 => n4201, B2 => n19029, C1 => n1896, C2 => 
                           n19023, A => n6614, ZN => n6610);
   U2877 : OAI221_X1 port map( B1 => n19005, B2 => n6559, C1 => n2119, C2 => 
                           n18999, A => n6615, ZN => n6609);
   U2878 : NOR4_X1 port map( A1 => n6543, A2 => n6544, A3 => n6545, A4 => n6546
                           , ZN => n6542);
   U2879 : OAI222_X1 port map( A1 => n1754, A2 => n19071, B1 => n3794, B2 => 
                           n19065, C1 => n3728, C2 => n19059, ZN => n6546);
   U2880 : OAI221_X1 port map( B1 => n4200, B2 => n19029, C1 => n1895, C2 => 
                           n19023, A => n6548, ZN => n6544);
   U2881 : OAI221_X1 port map( B1 => n19005, B2 => n6493, C1 => n2118, C2 => 
                           n18999, A => n6549, ZN => n6543);
   U2882 : NOR4_X1 port map( A1 => n6477, A2 => n6478, A3 => n6479, A4 => n6480
                           , ZN => n6476);
   U2883 : OAI222_X1 port map( A1 => n1753, A2 => n19071, B1 => n3793, B2 => 
                           n19065, C1 => n3727, C2 => n19059, ZN => n6480);
   U2884 : OAI221_X1 port map( B1 => n4199, B2 => n19029, C1 => n1894, C2 => 
                           n19023, A => n6482, ZN => n6478);
   U2885 : OAI221_X1 port map( B1 => n19005, B2 => n6427, C1 => n2117, C2 => 
                           n18999, A => n6483, ZN => n6477);
   U2886 : NOR4_X1 port map( A1 => n6411, A2 => n6412, A3 => n6413, A4 => n6414
                           , ZN => n6410);
   U2887 : OAI222_X1 port map( A1 => n1752, A2 => n19071, B1 => n3792, B2 => 
                           n19065, C1 => n3726, C2 => n19059, ZN => n6414);
   U2888 : OAI221_X1 port map( B1 => n4198, B2 => n19029, C1 => n1893, C2 => 
                           n19023, A => n6416, ZN => n6412);
   U2889 : OAI221_X1 port map( B1 => n19005, B2 => n6361, C1 => n2116, C2 => 
                           n18999, A => n6417, ZN => n6411);
   U2890 : NOR4_X1 port map( A1 => n6345, A2 => n6346, A3 => n6347, A4 => n6348
                           , ZN => n6344);
   U2891 : OAI222_X1 port map( A1 => n1751, A2 => n19071, B1 => n3791, B2 => 
                           n19065, C1 => n3725, C2 => n19059, ZN => n6348);
   U2892 : OAI221_X1 port map( B1 => n4197, B2 => n19029, C1 => n1892, C2 => 
                           n19023, A => n6350, ZN => n6346);
   U2893 : OAI221_X1 port map( B1 => n19005, B2 => n6295, C1 => n2115, C2 => 
                           n18999, A => n6351, ZN => n6345);
   U2894 : NOR4_X1 port map( A1 => n6279, A2 => n6280, A3 => n6281, A4 => n6282
                           , ZN => n6278);
   U2895 : OAI222_X1 port map( A1 => n1750, A2 => n19071, B1 => n3790, B2 => 
                           n19065, C1 => n3724, C2 => n19059, ZN => n6282);
   U2896 : OAI221_X1 port map( B1 => n4196, B2 => n19029, C1 => n1891, C2 => 
                           n19023, A => n6284, ZN => n6280);
   U2897 : OAI221_X1 port map( B1 => n19005, B2 => n6229, C1 => n2114, C2 => 
                           n18999, A => n6285, ZN => n6279);
   U2898 : NOR4_X1 port map( A1 => n6213, A2 => n6214, A3 => n6215, A4 => n6216
                           , ZN => n6212);
   U2899 : OAI222_X1 port map( A1 => n1749, A2 => n19071, B1 => n3789, B2 => 
                           n19065, C1 => n3723, C2 => n19059, ZN => n6216);
   U2900 : OAI221_X1 port map( B1 => n4195, B2 => n19029, C1 => n1890, C2 => 
                           n19023, A => n6218, ZN => n6214);
   U2901 : OAI221_X1 port map( B1 => n19005, B2 => n6163, C1 => n2113, C2 => 
                           n18999, A => n6219, ZN => n6213);
   U2902 : NOR4_X1 port map( A1 => n6147, A2 => n6148, A3 => n6149, A4 => n6150
                           , ZN => n6146);
   U2903 : OAI222_X1 port map( A1 => n1745, A2 => n19072, B1 => n3788, B2 => 
                           n19066, C1 => n3722, C2 => n19060, ZN => n6150);
   U2904 : OAI221_X1 port map( B1 => n4194, B2 => n19030, C1 => n1889, C2 => 
                           n19024, A => n6152, ZN => n6148);
   U2905 : OAI221_X1 port map( B1 => n19006, B2 => n6097, C1 => n2112, C2 => 
                           n19000, A => n6153, ZN => n6147);
   U2906 : NOR4_X1 port map( A1 => n6081, A2 => n6082, A3 => n6083, A4 => n6084
                           , ZN => n6080);
   U2907 : OAI222_X1 port map( A1 => n1744, A2 => n19072, B1 => n3787, B2 => 
                           n19066, C1 => n3721, C2 => n19060, ZN => n6084);
   U2908 : OAI221_X1 port map( B1 => n4193, B2 => n19030, C1 => n1888, C2 => 
                           n19024, A => n6086, ZN => n6082);
   U2909 : OAI221_X1 port map( B1 => n19006, B2 => n6029, C1 => n2111, C2 => 
                           n19000, A => n6087, ZN => n6081);
   U2910 : NOR4_X1 port map( A1 => n6013, A2 => n6014, A3 => n6015, A4 => n6016
                           , ZN => n6012);
   U2911 : OAI222_X1 port map( A1 => n1743, A2 => n19072, B1 => n3786, B2 => 
                           n19066, C1 => n3720, C2 => n19060, ZN => n6016);
   U2912 : OAI221_X1 port map( B1 => n4192, B2 => n19030, C1 => n1887, C2 => 
                           n19024, A => n6018, ZN => n6014);
   U2913 : OAI221_X1 port map( B1 => n19006, B2 => n5961, C1 => n2110, C2 => 
                           n19000, A => n6019, ZN => n6013);
   U2914 : NOR4_X1 port map( A1 => n5945, A2 => n5946, A3 => n5947, A4 => n5948
                           , ZN => n5944);
   U2915 : OAI222_X1 port map( A1 => n1742, A2 => n19072, B1 => n3785, B2 => 
                           n19066, C1 => n3719, C2 => n19060, ZN => n5948);
   U2916 : OAI221_X1 port map( B1 => n4191, B2 => n19030, C1 => n1886, C2 => 
                           n19024, A => n5950, ZN => n5946);
   U2917 : OAI221_X1 port map( B1 => n19006, B2 => n5894, C1 => n2109, C2 => 
                           n19000, A => n5951, ZN => n5945);
   U2918 : NOR4_X1 port map( A1 => n5878, A2 => n5879, A3 => n5880, A4 => n5881
                           , ZN => n5877);
   U2919 : OAI222_X1 port map( A1 => n1741, A2 => n19072, B1 => n3784, B2 => 
                           n19066, C1 => n3718, C2 => n19060, ZN => n5881);
   U2920 : OAI221_X1 port map( B1 => n4190, B2 => n19030, C1 => n1885, C2 => 
                           n19024, A => n5883, ZN => n5879);
   U2921 : OAI221_X1 port map( B1 => n19006, B2 => n5827, C1 => n2108, C2 => 
                           n19000, A => n5884, ZN => n5878);
   U2922 : NOR4_X1 port map( A1 => n5811, A2 => n5812, A3 => n5813, A4 => n5814
                           , ZN => n5810);
   U2923 : OAI222_X1 port map( A1 => n1740, A2 => n19072, B1 => n3783, B2 => 
                           n19066, C1 => n3717, C2 => n19060, ZN => n5814);
   U2924 : OAI221_X1 port map( B1 => n4189, B2 => n19030, C1 => n1884, C2 => 
                           n19024, A => n5816, ZN => n5812);
   U2925 : OAI221_X1 port map( B1 => n19006, B2 => n5755, C1 => n2107, C2 => 
                           n19000, A => n5817, ZN => n5811);
   U2926 : NOR4_X1 port map( A1 => n5739, A2 => n5740, A3 => n5741, A4 => n5742
                           , ZN => n5738);
   U2927 : OAI222_X1 port map( A1 => n1739, A2 => n19072, B1 => n3782, B2 => 
                           n19066, C1 => n3716, C2 => n19060, ZN => n5742);
   U2928 : OAI221_X1 port map( B1 => n4188, B2 => n19030, C1 => n1883, C2 => 
                           n19024, A => n5744, ZN => n5740);
   U2929 : OAI221_X1 port map( B1 => n19006, B2 => n5685, C1 => n2106, C2 => 
                           n19000, A => n5745, ZN => n5739);
   U2930 : NOR4_X1 port map( A1 => n5669, A2 => n5670, A3 => n5671, A4 => n5672
                           , ZN => n5668);
   U2931 : OAI222_X1 port map( A1 => n1738, A2 => n19072, B1 => n3781, B2 => 
                           n19066, C1 => n3715, C2 => n19060, ZN => n5672);
   U2932 : OAI221_X1 port map( B1 => n4187, B2 => n19030, C1 => n1882, C2 => 
                           n19024, A => n5674, ZN => n5670);
   U2933 : OAI221_X1 port map( B1 => n19006, B2 => n5617, C1 => n2105, C2 => 
                           n19000, A => n5675, ZN => n5669);
   U2934 : NOR4_X1 port map( A1 => n5601, A2 => n5602, A3 => n5603, A4 => n5604
                           , ZN => n5600);
   U2935 : OAI222_X1 port map( A1 => n1737, A2 => n19072, B1 => n3780, B2 => 
                           n19066, C1 => n3714, C2 => n19060, ZN => n5604);
   U2936 : OAI221_X1 port map( B1 => n4186, B2 => n19030, C1 => n1881, C2 => 
                           n19024, A => n5606, ZN => n5602);
   U2937 : OAI221_X1 port map( B1 => n19006, B2 => n5548, C1 => n2104, C2 => 
                           n19000, A => n5607, ZN => n5601);
   U2938 : NOR4_X1 port map( A1 => n5532, A2 => n5533, A3 => n5534, A4 => n5535
                           , ZN => n5531);
   U2939 : OAI222_X1 port map( A1 => n1736, A2 => n19072, B1 => n3779, B2 => 
                           n19066, C1 => n3713, C2 => n19060, ZN => n5535);
   U2940 : OAI221_X1 port map( B1 => n4185, B2 => n19030, C1 => n1880, C2 => 
                           n19024, A => n5537, ZN => n5533);
   U2941 : OAI221_X1 port map( B1 => n19006, B2 => n5479, C1 => n2103, C2 => 
                           n19000, A => n5538, ZN => n5532);
   U2942 : NOR4_X1 port map( A1 => n5463, A2 => n5464, A3 => n5465, A4 => n5466
                           , ZN => n5462);
   U2943 : OAI222_X1 port map( A1 => n1735, A2 => n19072, B1 => n3778, B2 => 
                           n19066, C1 => n3712, C2 => n19060, ZN => n5466);
   U2944 : OAI221_X1 port map( B1 => n4184, B2 => n19030, C1 => n1879, C2 => 
                           n19024, A => n5468, ZN => n5464);
   U2945 : OAI221_X1 port map( B1 => n19006, B2 => n5411, C1 => n2102, C2 => 
                           n19000, A => n5469, ZN => n5463);
   U2946 : NOR4_X1 port map( A1 => n5395, A2 => n5396, A3 => n5397, A4 => n5398
                           , ZN => n5394);
   U2947 : OAI222_X1 port map( A1 => n1734, A2 => n19072, B1 => n3777, B2 => 
                           n19066, C1 => n3711, C2 => n19060, ZN => n5398);
   U2948 : OAI221_X1 port map( B1 => n4183, B2 => n19030, C1 => n1878, C2 => 
                           n19024, A => n5400, ZN => n5396);
   U2949 : OAI221_X1 port map( B1 => n19006, B2 => n5341, C1 => n2101, C2 => 
                           n19000, A => n5401, ZN => n5395);
   U2950 : NOR4_X1 port map( A1 => n11666, A2 => n11667, A3 => n11668, A4 => 
                           n11669, ZN => n11665);
   U2951 : OAI222_X1 port map( A1 => n1796, A2 => n19068, B1 => n3836, B2 => 
                           n19062, C1 => n3770, C2 => n19056, ZN => n11669);
   U2952 : OAI221_X1 port map( B1 => n4242, B2 => n19026, C1 => n1937, C2 => 
                           n19020, A => n11685, ZN => n11667);
   U2953 : OAI221_X1 port map( B1 => n19002, B2 => n11555, C1 => n2192, C2 => 
                           n18996, A => n11689, ZN => n11666);
   U2954 : NOR4_X1 port map( A1 => n11538, A2 => n11539, A3 => n11540, A4 => 
                           n11541, ZN => n11537);
   U2955 : OAI222_X1 port map( A1 => n1795, A2 => n19068, B1 => n3835, B2 => 
                           n19062, C1 => n3769, C2 => n19056, ZN => n11541);
   U2956 : OAI221_X1 port map( B1 => n4241, B2 => n19026, C1 => n1936, C2 => 
                           n19020, A => n11544, ZN => n11539);
   U2957 : OAI221_X1 port map( B1 => n19002, B2 => n11487, C1 => n2189, C2 => 
                           n18996, A => n11545, ZN => n11538);
   U2958 : NOR4_X1 port map( A1 => n11471, A2 => n11472, A3 => n11473, A4 => 
                           n11474, ZN => n11470);
   U2959 : OAI222_X1 port map( A1 => n1794, A2 => n19068, B1 => n3834, B2 => 
                           n19062, C1 => n3768, C2 => n19056, ZN => n11474);
   U2960 : OAI221_X1 port map( B1 => n4240, B2 => n19026, C1 => n1935, C2 => 
                           n19020, A => n11476, ZN => n11472);
   U2961 : OAI221_X1 port map( B1 => n19002, B2 => n11420, C1 => n2186, C2 => 
                           n18996, A => n11477, ZN => n11471);
   U2962 : NOR4_X1 port map( A1 => n11404, A2 => n11405, A3 => n11406, A4 => 
                           n11407, ZN => n11403);
   U2963 : OAI222_X1 port map( A1 => n1793, A2 => n19068, B1 => n3833, B2 => 
                           n19062, C1 => n3767, C2 => n19056, ZN => n11407);
   U2964 : OAI221_X1 port map( B1 => n4239, B2 => n19026, C1 => n1934, C2 => 
                           n19020, A => n11409, ZN => n11405);
   U2965 : OAI221_X1 port map( B1 => n19002, B2 => n11353, C1 => n2183, C2 => 
                           n18996, A => n11410, ZN => n11404);
   U2966 : NOR4_X1 port map( A1 => n11337, A2 => n11338, A3 => n11339, A4 => 
                           n11340, ZN => n11336);
   U2967 : OAI222_X1 port map( A1 => n1792, A2 => n19068, B1 => n3832, B2 => 
                           n19062, C1 => n3766, C2 => n19056, ZN => n11340);
   U2968 : OAI221_X1 port map( B1 => n4238, B2 => n19026, C1 => n1933, C2 => 
                           n19020, A => n11342, ZN => n11338);
   U2969 : OAI221_X1 port map( B1 => n19002, B2 => n11286, C1 => n2180, C2 => 
                           n18996, A => n11343, ZN => n11337);
   U2970 : NOR4_X1 port map( A1 => n11269, A2 => n11270, A3 => n11271, A4 => 
                           n11272, ZN => n11268);
   U2971 : OAI222_X1 port map( A1 => n1791, A2 => n19068, B1 => n3831, B2 => 
                           n19062, C1 => n3765, C2 => n19056, ZN => n11272);
   U2972 : OAI221_X1 port map( B1 => n4237, B2 => n19026, C1 => n1932, C2 => 
                           n19020, A => n11274, ZN => n11270);
   U2973 : OAI221_X1 port map( B1 => n19002, B2 => n11218, C1 => n2177, C2 => 
                           n18996, A => n11275, ZN => n11269);
   U2974 : NOR4_X1 port map( A1 => n11202, A2 => n11203, A3 => n11204, A4 => 
                           n11205, ZN => n11201);
   U2975 : OAI222_X1 port map( A1 => n1790, A2 => n19068, B1 => n3830, B2 => 
                           n19062, C1 => n3764, C2 => n19056, ZN => n11205);
   U2976 : OAI221_X1 port map( B1 => n4236, B2 => n19026, C1 => n1931, C2 => 
                           n19020, A => n11207, ZN => n11203);
   U2977 : OAI221_X1 port map( B1 => n19002, B2 => n11151, C1 => n2174, C2 => 
                           n18996, A => n11208, ZN => n11202);
   U2978 : NOR4_X1 port map( A1 => n11135, A2 => n11136, A3 => n11137, A4 => 
                           n11138, ZN => n11134);
   U2979 : OAI222_X1 port map( A1 => n1789, A2 => n19068, B1 => n3829, B2 => 
                           n19062, C1 => n3763, C2 => n19056, ZN => n11138);
   U2980 : OAI221_X1 port map( B1 => n4235, B2 => n19026, C1 => n1930, C2 => 
                           n19020, A => n11140, ZN => n11136);
   U2981 : OAI221_X1 port map( B1 => n19002, B2 => n11084, C1 => n2171, C2 => 
                           n18996, A => n11141, ZN => n11135);
   U2982 : NOR4_X1 port map( A1 => n11068, A2 => n11069, A3 => n11070, A4 => 
                           n11071, ZN => n11067);
   U2983 : OAI222_X1 port map( A1 => n1788, A2 => n19068, B1 => n3828, B2 => 
                           n19062, C1 => n3762, C2 => n19056, ZN => n11071);
   U2984 : OAI221_X1 port map( B1 => n4234, B2 => n19026, C1 => n1929, C2 => 
                           n19020, A => n11073, ZN => n11069);
   U2985 : OAI221_X1 port map( B1 => n19002, B2 => n11017, C1 => n2168, C2 => 
                           n18996, A => n11074, ZN => n11068);
   U2986 : NOR4_X1 port map( A1 => n11000, A2 => n11001, A3 => n11002, A4 => 
                           n11003, ZN => n10999);
   U2987 : OAI222_X1 port map( A1 => n1787, A2 => n19068, B1 => n3827, B2 => 
                           n19062, C1 => n3761, C2 => n19056, ZN => n11003);
   U2988 : OAI221_X1 port map( B1 => n4233, B2 => n19026, C1 => n1928, C2 => 
                           n19020, A => n11005, ZN => n11001);
   U2989 : OAI221_X1 port map( B1 => n19002, B2 => n10949, C1 => n2165, C2 => 
                           n18996, A => n11006, ZN => n11000);
   U2990 : NOR4_X1 port map( A1 => n10933, A2 => n10934, A3 => n10935, A4 => 
                           n10936, ZN => n10932);
   U2991 : OAI222_X1 port map( A1 => n1786, A2 => n19068, B1 => n3826, B2 => 
                           n19062, C1 => n3760, C2 => n19056, ZN => n10936);
   U2992 : OAI221_X1 port map( B1 => n4232, B2 => n19026, C1 => n1927, C2 => 
                           n19020, A => n10938, ZN => n10934);
   U2993 : OAI221_X1 port map( B1 => n19002, B2 => n10882, C1 => n2162, C2 => 
                           n18996, A => n10939, ZN => n10933);
   U2994 : NOR4_X1 port map( A1 => n10866, A2 => n10867, A3 => n10868, A4 => 
                           n10869, ZN => n10865);
   U2995 : OAI222_X1 port map( A1 => n1785, A2 => n19068, B1 => n3825, B2 => 
                           n19062, C1 => n3759, C2 => n19056, ZN => n10869);
   U2996 : OAI221_X1 port map( B1 => n4231, B2 => n19026, C1 => n1926, C2 => 
                           n19020, A => n10871, ZN => n10867);
   U2997 : OAI221_X1 port map( B1 => n19002, B2 => n10815, C1 => n2159, C2 => 
                           n18996, A => n10872, ZN => n10866);
   U2998 : NOR4_X1 port map( A1 => n10798, A2 => n10799, A3 => n10800, A4 => 
                           n10802, ZN => n10797);
   U2999 : OAI222_X1 port map( A1 => n1784, A2 => n19069, B1 => n3824, B2 => 
                           n19063, C1 => n3758, C2 => n19057, ZN => n10802);
   U3000 : OAI221_X1 port map( B1 => n4230, B2 => n19027, C1 => n1925, C2 => 
                           n19021, A => n10804, ZN => n10799);
   U3001 : OAI221_X1 port map( B1 => n19003, B2 => n10747, C1 => n2156, C2 => 
                           n18997, A => n10805, ZN => n10798);
   U3002 : NOR4_X1 port map( A1 => n10731, A2 => n10732, A3 => n10733, A4 => 
                           n10734, ZN => n10730);
   U3003 : OAI222_X1 port map( A1 => n1783, A2 => n19069, B1 => n3823, B2 => 
                           n19063, C1 => n3757, C2 => n19057, ZN => n10734);
   U3004 : OAI221_X1 port map( B1 => n4229, B2 => n19027, C1 => n1924, C2 => 
                           n19021, A => n10736, ZN => n10732);
   U3005 : OAI221_X1 port map( B1 => n19003, B2 => n10680, C1 => n2153, C2 => 
                           n18997, A => n10737, ZN => n10731);
   U3006 : NOR4_X1 port map( A1 => n10664, A2 => n10665, A3 => n10666, A4 => 
                           n10667, ZN => n10663);
   U3007 : OAI222_X1 port map( A1 => n1782, A2 => n19069, B1 => n3822, B2 => 
                           n19063, C1 => n3756, C2 => n19057, ZN => n10667);
   U3008 : OAI221_X1 port map( B1 => n4228, B2 => n19027, C1 => n1923, C2 => 
                           n19021, A => n10669, ZN => n10665);
   U3009 : OAI221_X1 port map( B1 => n19003, B2 => n10613, C1 => n2150, C2 => 
                           n18997, A => n10670, ZN => n10664);
   U3010 : NOR4_X1 port map( A1 => n10597, A2 => n10598, A3 => n10599, A4 => 
                           n10600, ZN => n10596);
   U3011 : OAI222_X1 port map( A1 => n1781, A2 => n19069, B1 => n3821, B2 => 
                           n19063, C1 => n3755, C2 => n19057, ZN => n10600);
   U3012 : OAI221_X1 port map( B1 => n4227, B2 => n19027, C1 => n1922, C2 => 
                           n19021, A => n10602, ZN => n10598);
   U3013 : OAI221_X1 port map( B1 => n19003, B2 => n10546, C1 => n2147, C2 => 
                           n18997, A => n10603, ZN => n10597);
   U3014 : NOR4_X1 port map( A1 => n10529, A2 => n10530, A3 => n10531, A4 => 
                           n10532, ZN => n10528);
   U3015 : OAI222_X1 port map( A1 => n1780, A2 => n19069, B1 => n3820, B2 => 
                           n19063, C1 => n3754, C2 => n19057, ZN => n10532);
   U3016 : OAI221_X1 port map( B1 => n4226, B2 => n19027, C1 => n1921, C2 => 
                           n19021, A => n10534, ZN => n10530);
   U3017 : OAI221_X1 port map( B1 => n19003, B2 => n10478, C1 => n2144, C2 => 
                           n18997, A => n10535, ZN => n10529);
   U3018 : NOR4_X1 port map( A1 => n10462, A2 => n10463, A3 => n10464, A4 => 
                           n10465, ZN => n10461);
   U3019 : OAI222_X1 port map( A1 => n1779, A2 => n19069, B1 => n3819, B2 => 
                           n19063, C1 => n3753, C2 => n19057, ZN => n10465);
   U3020 : OAI221_X1 port map( B1 => n4225, B2 => n19027, C1 => n1920, C2 => 
                           n19021, A => n10467, ZN => n10463);
   U3021 : OAI221_X1 port map( B1 => n19003, B2 => n10411, C1 => n2143, C2 => 
                           n18997, A => n10468, ZN => n10462);
   U3022 : NOR4_X1 port map( A1 => n10395, A2 => n10396, A3 => n10397, A4 => 
                           n10398, ZN => n10394);
   U3023 : OAI222_X1 port map( A1 => n1778, A2 => n19069, B1 => n3818, B2 => 
                           n19063, C1 => n3752, C2 => n19057, ZN => n10398);
   U3024 : OAI221_X1 port map( B1 => n4224, B2 => n19027, C1 => n1919, C2 => 
                           n19021, A => n10400, ZN => n10396);
   U3025 : OAI221_X1 port map( B1 => n19003, B2 => n10344, C1 => n2142, C2 => 
                           n18997, A => n10401, ZN => n10395);
   U3026 : NOR4_X1 port map( A1 => n10328, A2 => n10329, A3 => n10330, A4 => 
                           n10331, ZN => n10327);
   U3027 : OAI222_X1 port map( A1 => n1777, A2 => n19069, B1 => n3817, B2 => 
                           n19063, C1 => n3751, C2 => n19057, ZN => n10331);
   U3028 : OAI221_X1 port map( B1 => n4223, B2 => n19027, C1 => n1918, C2 => 
                           n19021, A => n10333, ZN => n10329);
   U3029 : OAI221_X1 port map( B1 => n19003, B2 => n10277, C1 => n2141, C2 => 
                           n18997, A => n10334, ZN => n10328);
   U3030 : NOR4_X1 port map( A1 => n10260, A2 => n10261, A3 => n10262, A4 => 
                           n10263, ZN => n10259);
   U3031 : OAI222_X1 port map( A1 => n1776, A2 => n19069, B1 => n3816, B2 => 
                           n19063, C1 => n3750, C2 => n19057, ZN => n10263);
   U3032 : OAI221_X1 port map( B1 => n4222, B2 => n19027, C1 => n1917, C2 => 
                           n19021, A => n10265, ZN => n10261);
   U3033 : OAI221_X1 port map( B1 => n19003, B2 => n10209, C1 => n2140, C2 => 
                           n18997, A => n10266, ZN => n10260);
   U3034 : NOR4_X1 port map( A1 => n10193, A2 => n10194, A3 => n10195, A4 => 
                           n10196, ZN => n10192);
   U3035 : OAI222_X1 port map( A1 => n1775, A2 => n19069, B1 => n3815, B2 => 
                           n19063, C1 => n3749, C2 => n19057, ZN => n10196);
   U3036 : OAI221_X1 port map( B1 => n4221, B2 => n19027, C1 => n1916, C2 => 
                           n19021, A => n10198, ZN => n10194);
   U3037 : OAI221_X1 port map( B1 => n19003, B2 => n10142, C1 => n2139, C2 => 
                           n18997, A => n10199, ZN => n10193);
   U3038 : NOR4_X1 port map( A1 => n10126, A2 => n10127, A3 => n10128, A4 => 
                           n10129, ZN => n10125);
   U3039 : OAI222_X1 port map( A1 => n1774, A2 => n19069, B1 => n3814, B2 => 
                           n19063, C1 => n3748, C2 => n19057, ZN => n10129);
   U3040 : OAI221_X1 port map( B1 => n4220, B2 => n19027, C1 => n1915, C2 => 
                           n19021, A => n10131, ZN => n10127);
   U3041 : OAI221_X1 port map( B1 => n19003, B2 => n10075, C1 => n2138, C2 => 
                           n18997, A => n10132, ZN => n10126);
   U3042 : NOR4_X1 port map( A1 => n10058, A2 => n10060, A3 => n10061, A4 => 
                           n10062, ZN => n10057);
   U3043 : OAI222_X1 port map( A1 => n1773, A2 => n19069, B1 => n3813, B2 => 
                           n19063, C1 => n3747, C2 => n19057, ZN => n10062);
   U3044 : OAI221_X1 port map( B1 => n4219, B2 => n19027, C1 => n1914, C2 => 
                           n19021, A => n10064, ZN => n10060);
   U3045 : OAI221_X1 port map( B1 => n19003, B2 => n10008, C1 => n2137, C2 => 
                           n18997, A => n10065, ZN => n10058);
   U3046 : NOR4_X1 port map( A1 => n9991, A2 => n9992, A3 => n9993, A4 => n9994
                           , ZN => n9990);
   U3047 : OAI222_X1 port map( A1 => n1772, A2 => n19070, B1 => n3812, B2 => 
                           n19064, C1 => n3746, C2 => n19058, ZN => n9994);
   U3048 : OAI221_X1 port map( B1 => n4218, B2 => n19028, C1 => n1913, C2 => 
                           n19022, A => n9996, ZN => n9992);
   U3049 : OAI221_X1 port map( B1 => n19004, B2 => n9940, C1 => n2136, C2 => 
                           n18998, A => n9997, ZN => n9991);
   U3050 : NOR4_X1 port map( A1 => n9924, A2 => n9925, A3 => n9926, A4 => n9927
                           , ZN => n9923);
   U3051 : OAI222_X1 port map( A1 => n1771, A2 => n19070, B1 => n3811, B2 => 
                           n19064, C1 => n3745, C2 => n19058, ZN => n9927);
   U3052 : OAI221_X1 port map( B1 => n4217, B2 => n19028, C1 => n1912, C2 => 
                           n19022, A => n9929, ZN => n9925);
   U3053 : OAI221_X1 port map( B1 => n19004, B2 => n9873, C1 => n2135, C2 => 
                           n18998, A => n9930, ZN => n9924);
   U3054 : NOR4_X1 port map( A1 => n9857, A2 => n9858, A3 => n9859, A4 => n9860
                           , ZN => n9856);
   U3055 : OAI222_X1 port map( A1 => n1770, A2 => n19070, B1 => n3810, B2 => 
                           n19064, C1 => n3744, C2 => n19058, ZN => n9860);
   U3056 : OAI221_X1 port map( B1 => n4216, B2 => n19028, C1 => n1911, C2 => 
                           n19022, A => n9862, ZN => n9858);
   U3057 : OAI221_X1 port map( B1 => n19004, B2 => n9806, C1 => n2134, C2 => 
                           n18998, A => n9863, ZN => n9857);
   U3058 : NOR4_X1 port map( A1 => n9789, A2 => n9790, A3 => n9791, A4 => n9792
                           , ZN => n9788);
   U3059 : OAI222_X1 port map( A1 => n1769, A2 => n19070, B1 => n3809, B2 => 
                           n19064, C1 => n3743, C2 => n19058, ZN => n9792);
   U3060 : OAI221_X1 port map( B1 => n4215, B2 => n19028, C1 => n1910, C2 => 
                           n19022, A => n9794, ZN => n9790);
   U3061 : OAI221_X1 port map( B1 => n19004, B2 => n9738, C1 => n2133, C2 => 
                           n18998, A => n9796, ZN => n9789);
   U3062 : NOR4_X1 port map( A1 => n9722, A2 => n9723, A3 => n9724, A4 => n9725
                           , ZN => n9721);
   U3063 : OAI222_X1 port map( A1 => n1768, A2 => n19070, B1 => n3808, B2 => 
                           n19064, C1 => n3742, C2 => n19058, ZN => n9725);
   U3064 : OAI221_X1 port map( B1 => n4214, B2 => n19028, C1 => n1909, C2 => 
                           n19022, A => n9727, ZN => n9723);
   U3065 : OAI221_X1 port map( B1 => n19004, B2 => n9671, C1 => n2132, C2 => 
                           n18998, A => n9728, ZN => n9722);
   U3066 : NOR4_X1 port map( A1 => n9655, A2 => n9656, A3 => n9657, A4 => n9658
                           , ZN => n9654);
   U3067 : OAI222_X1 port map( A1 => n1767, A2 => n19070, B1 => n3807, B2 => 
                           n19064, C1 => n3741, C2 => n19058, ZN => n9658);
   U3068 : OAI221_X1 port map( B1 => n4213, B2 => n19028, C1 => n1908, C2 => 
                           n19022, A => n9660, ZN => n9656);
   U3069 : OAI221_X1 port map( B1 => n19004, B2 => n9604, C1 => n2131, C2 => 
                           n18998, A => n9661, ZN => n9655);
   U3070 : NOR4_X1 port map( A1 => n9588, A2 => n9589, A3 => n9590, A4 => n9591
                           , ZN => n9587);
   U3071 : OAI222_X1 port map( A1 => n1766, A2 => n19070, B1 => n3806, B2 => 
                           n19064, C1 => n3740, C2 => n19058, ZN => n9591);
   U3072 : OAI221_X1 port map( B1 => n4212, B2 => n19028, C1 => n1907, C2 => 
                           n19022, A => n9593, ZN => n9589);
   U3073 : OAI221_X1 port map( B1 => n19004, B2 => n9537, C1 => n2130, C2 => 
                           n18998, A => n9594, ZN => n9588);
   U3074 : NOR4_X1 port map( A1 => n9520, A2 => n9521, A3 => n9522, A4 => n9523
                           , ZN => n9519);
   U3075 : OAI222_X1 port map( A1 => n1765, A2 => n19070, B1 => n3805, B2 => 
                           n19064, C1 => n3739, C2 => n19058, ZN => n9523);
   U3076 : OAI221_X1 port map( B1 => n4211, B2 => n19028, C1 => n1906, C2 => 
                           n19022, A => n9525, ZN => n9521);
   U3077 : OAI221_X1 port map( B1 => n19004, B2 => n9469, C1 => n2129, C2 => 
                           n18998, A => n9526, ZN => n9520);
   U3078 : NOR4_X1 port map( A1 => n9453, A2 => n9454, A3 => n9455, A4 => n9456
                           , ZN => n9452);
   U3079 : OAI222_X1 port map( A1 => n1764, A2 => n19070, B1 => n3804, B2 => 
                           n19064, C1 => n3738, C2 => n19058, ZN => n9456);
   U3080 : OAI221_X1 port map( B1 => n4210, B2 => n19028, C1 => n1905, C2 => 
                           n19022, A => n9458, ZN => n9454);
   U3081 : OAI221_X1 port map( B1 => n19004, B2 => n9402, C1 => n2128, C2 => 
                           n18998, A => n9459, ZN => n9453);
   U3082 : NOR4_X1 port map( A1 => n9386, A2 => n9387, A3 => n9388, A4 => n9389
                           , ZN => n9385);
   U3083 : OAI222_X1 port map( A1 => n1763, A2 => n19070, B1 => n3803, B2 => 
                           n19064, C1 => n3737, C2 => n19058, ZN => n9389);
   U3084 : OAI221_X1 port map( B1 => n4209, B2 => n19028, C1 => n1904, C2 => 
                           n19022, A => n9391, ZN => n9387);
   U3085 : OAI221_X1 port map( B1 => n19004, B2 => n9335, C1 => n2127, C2 => 
                           n18998, A => n9392, ZN => n9386);
   U3086 : NOR4_X1 port map( A1 => n9319, A2 => n9320, A3 => n9321, A4 => n9322
                           , ZN => n9317);
   U3087 : OAI222_X1 port map( A1 => n1762, A2 => n19070, B1 => n3802, B2 => 
                           n19064, C1 => n3736, C2 => n19058, ZN => n9322);
   U3088 : OAI221_X1 port map( B1 => n4208, B2 => n19028, C1 => n1903, C2 => 
                           n19022, A => n9324, ZN => n9320);
   U3089 : OAI221_X1 port map( B1 => n19004, B2 => n9268, C1 => n2126, C2 => 
                           n18998, A => n9325, ZN => n9319);
   U3090 : NOR4_X1 port map( A1 => n7011, A2 => n7012, A3 => n7013, A4 => n7014
                           , ZN => n7010);
   U3091 : OAI222_X1 port map( A1 => n1761, A2 => n19070, B1 => n3801, B2 => 
                           n19064, C1 => n3735, C2 => n19058, ZN => n7014);
   U3092 : OAI221_X1 port map( B1 => n4207, B2 => n19028, C1 => n1902, C2 => 
                           n19022, A => n7016, ZN => n7012);
   U3093 : OAI221_X1 port map( B1 => n19004, B2 => n6961, C1 => n2125, C2 => 
                           n18998, A => n7017, ZN => n7011);
   U3094 : NOR4_X1 port map( A1 => n6944, A2 => n6945, A3 => n6947, A4 => n6948
                           , ZN => n6943);
   U3095 : OAI222_X1 port map( A1 => n1760, A2 => n19071, B1 => n3800, B2 => 
                           n19065, C1 => n3734, C2 => n19059, ZN => n6948);
   U3096 : OAI221_X1 port map( B1 => n4206, B2 => n19029, C1 => n1901, C2 => 
                           n19023, A => n6950, ZN => n6945);
   U3097 : OAI221_X1 port map( B1 => n19005, B2 => n6894, C1 => n2124, C2 => 
                           n18999, A => n6951, ZN => n6944);
   U3098 : NOR4_X1 port map( A1 => n6878, A2 => n6879, A3 => n6880, A4 => n6881
                           , ZN => n6877);
   U3099 : OAI222_X1 port map( A1 => n1759, A2 => n19071, B1 => n3799, B2 => 
                           n19065, C1 => n3733, C2 => n19059, ZN => n6881);
   U3100 : OAI221_X1 port map( B1 => n4205, B2 => n19029, C1 => n1900, C2 => 
                           n19023, A => n6883, ZN => n6879);
   U3101 : OAI221_X1 port map( B1 => n19005, B2 => n6827, C1 => n2123, C2 => 
                           n18999, A => n6884, ZN => n6878);
   U3102 : NOR4_X1 port map( A1 => n11628, A2 => n11629, A3 => n11630, A4 => 
                           n11631, ZN => n11627);
   U3103 : OAI221_X1 port map( B1 => n1937, B2 => n19267, C1 => n19266, C2 => 
                           n2145, A => n11632, ZN => n11631);
   U3104 : OAI221_X1 port map( B1 => n4921, B2 => n19243, C1 => n2441, C2 => 
                           n19237, A => n11638, ZN => n11630);
   U3105 : OAI221_X1 port map( B1 => n1863, B2 => n19195, C1 => n4242, C2 => 
                           n19189, A => n11646, ZN => n11628);
   U3106 : NOR4_X1 port map( A1 => n11580, A2 => n11581, A3 => n11582, A4 => 
                           n11583, ZN => n11579);
   U3107 : OAI221_X1 port map( B1 => n1863, B2 => n19394, C1 => n4242, C2 => 
                           n19388, A => n11604, ZN => n11580);
   U3108 : OAI221_X1 port map( B1 => n1937, B2 => n19466, C1 => n19465, C2 => 
                           n2146, A => n11584, ZN => n11583);
   U3109 : OAI221_X1 port map( B1 => n3366, B2 => n19418, C1 => n4850, C2 => 
                           n19412, A => n11597, ZN => n11581);
   U3110 : NOR4_X1 port map( A1 => n11520, A2 => n11521, A3 => n11522, A4 => 
                           n11523, ZN => n11519);
   U3111 : OAI221_X1 port map( B1 => n1936, B2 => n19267, C1 => n19266, C2 => 
                           n2148, A => n11524, ZN => n11523);
   U3112 : OAI221_X1 port map( B1 => n4920, B2 => n19243, C1 => n2440, C2 => 
                           n19237, A => n11525, ZN => n11522);
   U3113 : OAI221_X1 port map( B1 => n1862, B2 => n19195, C1 => n4241, C2 => 
                           n19189, A => n11527, ZN => n11520);
   U3114 : NOR4_X1 port map( A1 => n11493, A2 => n11494, A3 => n11495, A4 => 
                           n11496, ZN => n11492);
   U3115 : OAI221_X1 port map( B1 => n1862, B2 => n19394, C1 => n4241, C2 => 
                           n19388, A => n11505, ZN => n11493);
   U3116 : OAI221_X1 port map( B1 => n1936, B2 => n19466, C1 => n19465, C2 => 
                           n2149, A => n11497, ZN => n11496);
   U3117 : OAI221_X1 port map( B1 => n3365, B2 => n19418, C1 => n4849, C2 => 
                           n19412, A => n11502, ZN => n11494);
   U3118 : NOR4_X1 port map( A1 => n11453, A2 => n11454, A3 => n11455, A4 => 
                           n11456, ZN => n11452);
   U3119 : OAI221_X1 port map( B1 => n1935, B2 => n19267, C1 => n19266, C2 => 
                           n2151, A => n11457, ZN => n11456);
   U3120 : OAI221_X1 port map( B1 => n4919, B2 => n19243, C1 => n2439, C2 => 
                           n19237, A => n11458, ZN => n11455);
   U3121 : OAI221_X1 port map( B1 => n1861, B2 => n19195, C1 => n4240, C2 => 
                           n19189, A => n11460, ZN => n11453);
   U3122 : NOR4_X1 port map( A1 => n11425, A2 => n11426, A3 => n11427, A4 => 
                           n11428, ZN => n11424);
   U3123 : OAI221_X1 port map( B1 => n1861, B2 => n19394, C1 => n4240, C2 => 
                           n19388, A => n11438, ZN => n11425);
   U3124 : OAI221_X1 port map( B1 => n1935, B2 => n19466, C1 => n19465, C2 => 
                           n2152, A => n11429, ZN => n11428);
   U3125 : OAI221_X1 port map( B1 => n3364, B2 => n19418, C1 => n4848, C2 => 
                           n19412, A => n11434, ZN => n11426);
   U3126 : NOR4_X1 port map( A1 => n11386, A2 => n11387, A3 => n11388, A4 => 
                           n11389, ZN => n11385);
   U3127 : OAI221_X1 port map( B1 => n1934, B2 => n19267, C1 => n19266, C2 => 
                           n2154, A => n11390, ZN => n11389);
   U3128 : OAI221_X1 port map( B1 => n4918, B2 => n19243, C1 => n2438, C2 => 
                           n19237, A => n11391, ZN => n11388);
   U3129 : OAI221_X1 port map( B1 => n1860, B2 => n19195, C1 => n4239, C2 => 
                           n19189, A => n11393, ZN => n11386);
   U3130 : NOR4_X1 port map( A1 => n11358, A2 => n11359, A3 => n11360, A4 => 
                           n11361, ZN => n11357);
   U3131 : OAI221_X1 port map( B1 => n1860, B2 => n19394, C1 => n4239, C2 => 
                           n19388, A => n11370, ZN => n11358);
   U3132 : OAI221_X1 port map( B1 => n1934, B2 => n19466, C1 => n19465, C2 => 
                           n2155, A => n11362, ZN => n11361);
   U3133 : OAI221_X1 port map( B1 => n3363, B2 => n19418, C1 => n4847, C2 => 
                           n19412, A => n11367, ZN => n11359);
   U3134 : NOR4_X1 port map( A1 => n11318, A2 => n11319, A3 => n11320, A4 => 
                           n11321, ZN => n11317);
   U3135 : OAI221_X1 port map( B1 => n1933, B2 => n19267, C1 => n19265, C2 => 
                           n2157, A => n11322, ZN => n11321);
   U3136 : OAI221_X1 port map( B1 => n4917, B2 => n19243, C1 => n2437, C2 => 
                           n19237, A => n11323, ZN => n11320);
   U3137 : OAI221_X1 port map( B1 => n1859, B2 => n19195, C1 => n4238, C2 => 
                           n19189, A => n11325, ZN => n11318);
   U3138 : NOR4_X1 port map( A1 => n11291, A2 => n11292, A3 => n11293, A4 => 
                           n11294, ZN => n11290);
   U3139 : OAI221_X1 port map( B1 => n1859, B2 => n19394, C1 => n4238, C2 => 
                           n19388, A => n11303, ZN => n11291);
   U3140 : OAI221_X1 port map( B1 => n1933, B2 => n19466, C1 => n19464, C2 => 
                           n2158, A => n11295, ZN => n11294);
   U3141 : OAI221_X1 port map( B1 => n3362, B2 => n19418, C1 => n4846, C2 => 
                           n19412, A => n11300, ZN => n11292);
   U3142 : NOR4_X1 port map( A1 => n11251, A2 => n11252, A3 => n11253, A4 => 
                           n11254, ZN => n11250);
   U3143 : OAI221_X1 port map( B1 => n1932, B2 => n19267, C1 => n19265, C2 => 
                           n2160, A => n11255, ZN => n11254);
   U3144 : OAI221_X1 port map( B1 => n4916, B2 => n19243, C1 => n2436, C2 => 
                           n19237, A => n11256, ZN => n11253);
   U3145 : OAI221_X1 port map( B1 => n1858, B2 => n19195, C1 => n4237, C2 => 
                           n19189, A => n11258, ZN => n11251);
   U3146 : NOR4_X1 port map( A1 => n11223, A2 => n11224, A3 => n11226, A4 => 
                           n11227, ZN => n11222);
   U3147 : OAI221_X1 port map( B1 => n1858, B2 => n19394, C1 => n4237, C2 => 
                           n19388, A => n11236, ZN => n11223);
   U3148 : OAI221_X1 port map( B1 => n1932, B2 => n19466, C1 => n19464, C2 => 
                           n2161, A => n11228, ZN => n11227);
   U3149 : OAI221_X1 port map( B1 => n3361, B2 => n19418, C1 => n4845, C2 => 
                           n19412, A => n11233, ZN => n11224);
   U3150 : NOR4_X1 port map( A1 => n11184, A2 => n11185, A3 => n11186, A4 => 
                           n11187, ZN => n11183);
   U3151 : OAI221_X1 port map( B1 => n1931, B2 => n19267, C1 => n19265, C2 => 
                           n2163, A => n11188, ZN => n11187);
   U3152 : OAI221_X1 port map( B1 => n4915, B2 => n19243, C1 => n2435, C2 => 
                           n19237, A => n11189, ZN => n11186);
   U3153 : OAI221_X1 port map( B1 => n1857, B2 => n19195, C1 => n4236, C2 => 
                           n19189, A => n11191, ZN => n11184);
   U3154 : NOR4_X1 port map( A1 => n11156, A2 => n11157, A3 => n11158, A4 => 
                           n11159, ZN => n11155);
   U3155 : OAI221_X1 port map( B1 => n1857, B2 => n19394, C1 => n4236, C2 => 
                           n19388, A => n11168, ZN => n11156);
   U3156 : OAI221_X1 port map( B1 => n1931, B2 => n19466, C1 => n19464, C2 => 
                           n2164, A => n11160, ZN => n11159);
   U3157 : OAI221_X1 port map( B1 => n3360, B2 => n19418, C1 => n4844, C2 => 
                           n19412, A => n11165, ZN => n11157);
   U3158 : NOR4_X1 port map( A1 => n11116, A2 => n11117, A3 => n11118, A4 => 
                           n11120, ZN => n11115);
   U3159 : OAI221_X1 port map( B1 => n1930, B2 => n19267, C1 => n19265, C2 => 
                           n2166, A => n11121, ZN => n11120);
   U3160 : OAI221_X1 port map( B1 => n4914, B2 => n19243, C1 => n2434, C2 => 
                           n19237, A => n11122, ZN => n11118);
   U3161 : OAI221_X1 port map( B1 => n1856, B2 => n19195, C1 => n4235, C2 => 
                           n19189, A => n11124, ZN => n11116);
   U3162 : NOR4_X1 port map( A1 => n11089, A2 => n11090, A3 => n11091, A4 => 
                           n11092, ZN => n11088);
   U3163 : OAI221_X1 port map( B1 => n1856, B2 => n19394, C1 => n4235, C2 => 
                           n19388, A => n11101, ZN => n11089);
   U3164 : OAI221_X1 port map( B1 => n1930, B2 => n19466, C1 => n19464, C2 => 
                           n2167, A => n11093, ZN => n11092);
   U3165 : OAI221_X1 port map( B1 => n3359, B2 => n19418, C1 => n4843, C2 => 
                           n19412, A => n11098, ZN => n11090);
   U3166 : NOR4_X1 port map( A1 => n11049, A2 => n11050, A3 => n11051, A4 => 
                           n11052, ZN => n11048);
   U3167 : OAI221_X1 port map( B1 => n1929, B2 => n19267, C1 => n19265, C2 => 
                           n2169, A => n11053, ZN => n11052);
   U3168 : OAI221_X1 port map( B1 => n4913, B2 => n19243, C1 => n2433, C2 => 
                           n19237, A => n11054, ZN => n11051);
   U3169 : OAI221_X1 port map( B1 => n1855, B2 => n19195, C1 => n4234, C2 => 
                           n19189, A => n11056, ZN => n11049);
   U3170 : NOR4_X1 port map( A1 => n11022, A2 => n11023, A3 => n11024, A4 => 
                           n11025, ZN => n11021);
   U3171 : OAI221_X1 port map( B1 => n1855, B2 => n19394, C1 => n4234, C2 => 
                           n19388, A => n11034, ZN => n11022);
   U3172 : OAI221_X1 port map( B1 => n1929, B2 => n19466, C1 => n19464, C2 => 
                           n2170, A => n11026, ZN => n11025);
   U3173 : OAI221_X1 port map( B1 => n3358, B2 => n19418, C1 => n4842, C2 => 
                           n19412, A => n11031, ZN => n11023);
   U3174 : NOR4_X1 port map( A1 => n10982, A2 => n10983, A3 => n10984, A4 => 
                           n10985, ZN => n10981);
   U3175 : OAI221_X1 port map( B1 => n1928, B2 => n19267, C1 => n19265, C2 => 
                           n2172, A => n10986, ZN => n10985);
   U3176 : OAI221_X1 port map( B1 => n4912, B2 => n19243, C1 => n2432, C2 => 
                           n19237, A => n10987, ZN => n10984);
   U3177 : OAI221_X1 port map( B1 => n1854, B2 => n19195, C1 => n4233, C2 => 
                           n19189, A => n10989, ZN => n10982);
   U3178 : NOR4_X1 port map( A1 => n10954, A2 => n10955, A3 => n10956, A4 => 
                           n10957, ZN => n10953);
   U3179 : OAI221_X1 port map( B1 => n1854, B2 => n19394, C1 => n4233, C2 => 
                           n19388, A => n10967, ZN => n10954);
   U3180 : OAI221_X1 port map( B1 => n1928, B2 => n19466, C1 => n19464, C2 => 
                           n2173, A => n10958, ZN => n10957);
   U3181 : OAI221_X1 port map( B1 => n3357, B2 => n19418, C1 => n4841, C2 => 
                           n19412, A => n10964, ZN => n10955);
   U3182 : NOR4_X1 port map( A1 => n10915, A2 => n10916, A3 => n10917, A4 => 
                           n10918, ZN => n10914);
   U3183 : OAI221_X1 port map( B1 => n1927, B2 => n19267, C1 => n19265, C2 => 
                           n2175, A => n10919, ZN => n10918);
   U3184 : OAI221_X1 port map( B1 => n4911, B2 => n19243, C1 => n2431, C2 => 
                           n19237, A => n10920, ZN => n10917);
   U3185 : OAI221_X1 port map( B1 => n1853, B2 => n19195, C1 => n4232, C2 => 
                           n19189, A => n10922, ZN => n10915);
   U3186 : NOR4_X1 port map( A1 => n10887, A2 => n10888, A3 => n10889, A4 => 
                           n10890, ZN => n10886);
   U3187 : OAI221_X1 port map( B1 => n1853, B2 => n19394, C1 => n4232, C2 => 
                           n19388, A => n10899, ZN => n10887);
   U3188 : OAI221_X1 port map( B1 => n1927, B2 => n19466, C1 => n19464, C2 => 
                           n2176, A => n10891, ZN => n10890);
   U3189 : OAI221_X1 port map( B1 => n3356, B2 => n19418, C1 => n4840, C2 => 
                           n19412, A => n10896, ZN => n10888);
   U3190 : NOR4_X1 port map( A1 => n10847, A2 => n10848, A3 => n10849, A4 => 
                           n10850, ZN => n10846);
   U3191 : OAI221_X1 port map( B1 => n1926, B2 => n19267, C1 => n19265, C2 => 
                           n2178, A => n10851, ZN => n10850);
   U3192 : OAI221_X1 port map( B1 => n4910, B2 => n19243, C1 => n2430, C2 => 
                           n19237, A => n10852, ZN => n10849);
   U3193 : OAI221_X1 port map( B1 => n1852, B2 => n19195, C1 => n4231, C2 => 
                           n19189, A => n10855, ZN => n10847);
   U3194 : NOR4_X1 port map( A1 => n10820, A2 => n10821, A3 => n10822, A4 => 
                           n10823, ZN => n10819);
   U3195 : OAI221_X1 port map( B1 => n1852, B2 => n19394, C1 => n4231, C2 => 
                           n19388, A => n10832, ZN => n10820);
   U3196 : OAI221_X1 port map( B1 => n1926, B2 => n19466, C1 => n19464, C2 => 
                           n2179, A => n10824, ZN => n10823);
   U3197 : OAI221_X1 port map( B1 => n3355, B2 => n19418, C1 => n4839, C2 => 
                           n19412, A => n10829, ZN => n10821);
   U3198 : NOR4_X1 port map( A1 => n10780, A2 => n10781, A3 => n10782, A4 => 
                           n10783, ZN => n10779);
   U3199 : OAI221_X1 port map( B1 => n1925, B2 => n19268, C1 => n19265, C2 => 
                           n2181, A => n10784, ZN => n10783);
   U3200 : OAI221_X1 port map( B1 => n4909, B2 => n19244, C1 => n2429, C2 => 
                           n19238, A => n10785, ZN => n10782);
   U3201 : OAI221_X1 port map( B1 => n1851, B2 => n19196, C1 => n4230, C2 => 
                           n19190, A => n10787, ZN => n10780);
   U3202 : NOR4_X1 port map( A1 => n10753, A2 => n10754, A3 => n10755, A4 => 
                           n10756, ZN => n10752);
   U3203 : OAI221_X1 port map( B1 => n1851, B2 => n19395, C1 => n4230, C2 => 
                           n19389, A => n10765, ZN => n10753);
   U3204 : OAI221_X1 port map( B1 => n1925, B2 => n19467, C1 => n19464, C2 => 
                           n2182, A => n10757, ZN => n10756);
   U3205 : OAI221_X1 port map( B1 => n3354, B2 => n19419, C1 => n4838, C2 => 
                           n19413, A => n10762, ZN => n10754);
   U3206 : NOR4_X1 port map( A1 => n10713, A2 => n10714, A3 => n10715, A4 => 
                           n10716, ZN => n10712);
   U3207 : OAI221_X1 port map( B1 => n1924, B2 => n19268, C1 => n19265, C2 => 
                           n2184, A => n10717, ZN => n10716);
   U3208 : OAI221_X1 port map( B1 => n4908, B2 => n19244, C1 => n2428, C2 => 
                           n19238, A => n10718, ZN => n10715);
   U3209 : OAI221_X1 port map( B1 => n1850, B2 => n19196, C1 => n4229, C2 => 
                           n19190, A => n10720, ZN => n10713);
   U3210 : NOR4_X1 port map( A1 => n10685, A2 => n10686, A3 => n10687, A4 => 
                           n10688, ZN => n10684);
   U3211 : OAI221_X1 port map( B1 => n1850, B2 => n19395, C1 => n4229, C2 => 
                           n19389, A => n10698, ZN => n10685);
   U3212 : OAI221_X1 port map( B1 => n1924, B2 => n19467, C1 => n19464, C2 => 
                           n2185, A => n10689, ZN => n10688);
   U3213 : OAI221_X1 port map( B1 => n3353, B2 => n19419, C1 => n4837, C2 => 
                           n19413, A => n10694, ZN => n10686);
   U3214 : NOR4_X1 port map( A1 => n10646, A2 => n10647, A3 => n10648, A4 => 
                           n10649, ZN => n10645);
   U3215 : OAI221_X1 port map( B1 => n1923, B2 => n19268, C1 => n19265, C2 => 
                           n2187, A => n10650, ZN => n10649);
   U3216 : OAI221_X1 port map( B1 => n4907, B2 => n19244, C1 => n2427, C2 => 
                           n19238, A => n10651, ZN => n10648);
   U3217 : OAI221_X1 port map( B1 => n1849, B2 => n19196, C1 => n4228, C2 => 
                           n19190, A => n10653, ZN => n10646);
   U3218 : NOR4_X1 port map( A1 => n10618, A2 => n10619, A3 => n10620, A4 => 
                           n10621, ZN => n10617);
   U3219 : OAI221_X1 port map( B1 => n1849, B2 => n19395, C1 => n4228, C2 => 
                           n19389, A => n10630, ZN => n10618);
   U3220 : OAI221_X1 port map( B1 => n1923, B2 => n19467, C1 => n19464, C2 => 
                           n2188, A => n10622, ZN => n10621);
   U3221 : OAI221_X1 port map( B1 => n3352, B2 => n19419, C1 => n4836, C2 => 
                           n19413, A => n10627, ZN => n10619);
   U3222 : NOR4_X1 port map( A1 => n10578, A2 => n10579, A3 => n10580, A4 => 
                           n10581, ZN => n10577);
   U3223 : OAI221_X1 port map( B1 => n1922, B2 => n19268, C1 => n19265, C2 => 
                           n2190, A => n10582, ZN => n10581);
   U3224 : OAI221_X1 port map( B1 => n4906, B2 => n19244, C1 => n2426, C2 => 
                           n19238, A => n10583, ZN => n10580);
   U3225 : OAI221_X1 port map( B1 => n1848, B2 => n19196, C1 => n4227, C2 => 
                           n19190, A => n10585, ZN => n10578);
   U3226 : NOR4_X1 port map( A1 => n10551, A2 => n10552, A3 => n10553, A4 => 
                           n10554, ZN => n10550);
   U3227 : OAI221_X1 port map( B1 => n1848, B2 => n19395, C1 => n4227, C2 => 
                           n19389, A => n10563, ZN => n10551);
   U3228 : OAI221_X1 port map( B1 => n1922, B2 => n19467, C1 => n19464, C2 => 
                           n2191, A => n10555, ZN => n10554);
   U3229 : OAI221_X1 port map( B1 => n3351, B2 => n19419, C1 => n4835, C2 => 
                           n19413, A => n10560, ZN => n10552);
   U3230 : NOR4_X1 port map( A1 => n10511, A2 => n10512, A3 => n10513, A4 => 
                           n10514, ZN => n10510);
   U3231 : OAI221_X1 port map( B1 => n1921, B2 => n19268, C1 => n19264, C2 => 
                           n2193, A => n10515, ZN => n10514);
   U3232 : OAI221_X1 port map( B1 => n4905, B2 => n19244, C1 => n2425, C2 => 
                           n19238, A => n10516, ZN => n10513);
   U3233 : OAI221_X1 port map( B1 => n1847, B2 => n19196, C1 => n4226, C2 => 
                           n19190, A => n10518, ZN => n10511);
   U3234 : NOR4_X1 port map( A1 => n10484, A2 => n10485, A3 => n10486, A4 => 
                           n10487, ZN => n10482);
   U3235 : OAI221_X1 port map( B1 => n1847, B2 => n19395, C1 => n4226, C2 => 
                           n19389, A => n10496, ZN => n10484);
   U3236 : OAI221_X1 port map( B1 => n1921, B2 => n19467, C1 => n19463, C2 => 
                           n2194, A => n10488, ZN => n10487);
   U3237 : OAI221_X1 port map( B1 => n3350, B2 => n19419, C1 => n4834, C2 => 
                           n19413, A => n10493, ZN => n10485);
   U3238 : NOR4_X1 port map( A1 => n10444, A2 => n10445, A3 => n10446, A4 => 
                           n10447, ZN => n10443);
   U3239 : OAI221_X1 port map( B1 => n1920, B2 => n19268, C1 => n19264, C2 => 
                           n2196, A => n10448, ZN => n10447);
   U3240 : OAI221_X1 port map( B1 => n4904, B2 => n19244, C1 => n2424, C2 => 
                           n19238, A => n10449, ZN => n10446);
   U3241 : OAI221_X1 port map( B1 => n1846, B2 => n19196, C1 => n4225, C2 => 
                           n19190, A => n10451, ZN => n10444);
   U3242 : NOR4_X1 port map( A1 => n10416, A2 => n10417, A3 => n10418, A4 => 
                           n10419, ZN => n10415);
   U3243 : OAI221_X1 port map( B1 => n1846, B2 => n19395, C1 => n4225, C2 => 
                           n19389, A => n10428, ZN => n10416);
   U3244 : OAI221_X1 port map( B1 => n1920, B2 => n19467, C1 => n19463, C2 => 
                           n2197, A => n10420, ZN => n10419);
   U3245 : OAI221_X1 port map( B1 => n3349, B2 => n19419, C1 => n4833, C2 => 
                           n19413, A => n10425, ZN => n10417);
   U3246 : NOR4_X1 port map( A1 => n10376, A2 => n10378, A3 => n10379, A4 => 
                           n10380, ZN => n10375);
   U3247 : OAI221_X1 port map( B1 => n1919, B2 => n19268, C1 => n19264, C2 => 
                           n2199, A => n10381, ZN => n10380);
   U3248 : OAI221_X1 port map( B1 => n4903, B2 => n19244, C1 => n2423, C2 => 
                           n19238, A => n10382, ZN => n10379);
   U3249 : OAI221_X1 port map( B1 => n1845, B2 => n19196, C1 => n4224, C2 => 
                           n19190, A => n10384, ZN => n10376);
   U3250 : NOR4_X1 port map( A1 => n10349, A2 => n10350, A3 => n10351, A4 => 
                           n10352, ZN => n10348);
   U3251 : OAI221_X1 port map( B1 => n1845, B2 => n19395, C1 => n4224, C2 => 
                           n19389, A => n10361, ZN => n10349);
   U3252 : OAI221_X1 port map( B1 => n1919, B2 => n19467, C1 => n19463, C2 => 
                           n2200, A => n10353, ZN => n10352);
   U3253 : OAI221_X1 port map( B1 => n3348, B2 => n19419, C1 => n4832, C2 => 
                           n19413, A => n10358, ZN => n10350);
   U3254 : NOR4_X1 port map( A1 => n10309, A2 => n10310, A3 => n10311, A4 => 
                           n10312, ZN => n10308);
   U3255 : OAI221_X1 port map( B1 => n1918, B2 => n19268, C1 => n19264, C2 => 
                           n2202, A => n10313, ZN => n10312);
   U3256 : OAI221_X1 port map( B1 => n4902, B2 => n19244, C1 => n2422, C2 => 
                           n19238, A => n10314, ZN => n10311);
   U3257 : OAI221_X1 port map( B1 => n1844, B2 => n19196, C1 => n4223, C2 => 
                           n19190, A => n10316, ZN => n10309);
   U3258 : NOR4_X1 port map( A1 => n10282, A2 => n10283, A3 => n10284, A4 => 
                           n10285, ZN => n10281);
   U3259 : OAI221_X1 port map( B1 => n1844, B2 => n19395, C1 => n4223, C2 => 
                           n19389, A => n10294, ZN => n10282);
   U3260 : OAI221_X1 port map( B1 => n1918, B2 => n19467, C1 => n19463, C2 => 
                           n2203, A => n10286, ZN => n10285);
   U3261 : OAI221_X1 port map( B1 => n3347, B2 => n19419, C1 => n4831, C2 => 
                           n19413, A => n10291, ZN => n10283);
   U3262 : NOR4_X1 port map( A1 => n10242, A2 => n10243, A3 => n10244, A4 => 
                           n10245, ZN => n10241);
   U3263 : OAI221_X1 port map( B1 => n1917, B2 => n19268, C1 => n19264, C2 => 
                           n2205, A => n10246, ZN => n10245);
   U3264 : OAI221_X1 port map( B1 => n4901, B2 => n19244, C1 => n2421, C2 => 
                           n19238, A => n10247, ZN => n10244);
   U3265 : OAI221_X1 port map( B1 => n1843, B2 => n19196, C1 => n4222, C2 => 
                           n19190, A => n10249, ZN => n10242);
   U3266 : NOR4_X1 port map( A1 => n10214, A2 => n10215, A3 => n10216, A4 => 
                           n10217, ZN => n10213);
   U3267 : OAI221_X1 port map( B1 => n1843, B2 => n19395, C1 => n4222, C2 => 
                           n19389, A => n10227, ZN => n10214);
   U3268 : OAI221_X1 port map( B1 => n1917, B2 => n19467, C1 => n19463, C2 => 
                           n2206, A => n10219, ZN => n10217);
   U3269 : OAI221_X1 port map( B1 => n3346, B2 => n19419, C1 => n4830, C2 => 
                           n19413, A => n10224, ZN => n10215);
   U3270 : NOR4_X1 port map( A1 => n10175, A2 => n10176, A3 => n10177, A4 => 
                           n10178, ZN => n10174);
   U3271 : OAI221_X1 port map( B1 => n1916, B2 => n19268, C1 => n19264, C2 => 
                           n2208, A => n10179, ZN => n10178);
   U3272 : OAI221_X1 port map( B1 => n4900, B2 => n19244, C1 => n2420, C2 => 
                           n19238, A => n10180, ZN => n10177);
   U3273 : OAI221_X1 port map( B1 => n1842, B2 => n19196, C1 => n4221, C2 => 
                           n19190, A => n10182, ZN => n10175);
   U3274 : NOR4_X1 port map( A1 => n10147, A2 => n10148, A3 => n10149, A4 => 
                           n10150, ZN => n10146);
   U3275 : OAI221_X1 port map( B1 => n1842, B2 => n19395, C1 => n4221, C2 => 
                           n19389, A => n10159, ZN => n10147);
   U3276 : OAI221_X1 port map( B1 => n1916, B2 => n19467, C1 => n19463, C2 => 
                           n2209, A => n10151, ZN => n10150);
   U3277 : OAI221_X1 port map( B1 => n3345, B2 => n19419, C1 => n4829, C2 => 
                           n19413, A => n10156, ZN => n10148);
   U3278 : NOR4_X1 port map( A1 => n10107, A2 => n10108, A3 => n10109, A4 => 
                           n10110, ZN => n10106);
   U3279 : OAI221_X1 port map( B1 => n1915, B2 => n19268, C1 => n19264, C2 => 
                           n2211, A => n10111, ZN => n10110);
   U3280 : OAI221_X1 port map( B1 => n4899, B2 => n19244, C1 => n2419, C2 => 
                           n19238, A => n10113, ZN => n10109);
   U3281 : OAI221_X1 port map( B1 => n1841, B2 => n19196, C1 => n4220, C2 => 
                           n19190, A => n10115, ZN => n10107);
   U3282 : NOR4_X1 port map( A1 => n10080, A2 => n10081, A3 => n10082, A4 => 
                           n10083, ZN => n10079);
   U3283 : OAI221_X1 port map( B1 => n1841, B2 => n19395, C1 => n4220, C2 => 
                           n19389, A => n10092, ZN => n10080);
   U3284 : OAI221_X1 port map( B1 => n1915, B2 => n19467, C1 => n19463, C2 => 
                           n2212, A => n10084, ZN => n10083);
   U3285 : OAI221_X1 port map( B1 => n3344, B2 => n19419, C1 => n4828, C2 => 
                           n19413, A => n10089, ZN => n10081);
   U3286 : NOR4_X1 port map( A1 => n10040, A2 => n10041, A3 => n10042, A4 => 
                           n10043, ZN => n10039);
   U3287 : OAI221_X1 port map( B1 => n1914, B2 => n19268, C1 => n19264, C2 => 
                           n2214, A => n10044, ZN => n10043);
   U3288 : OAI221_X1 port map( B1 => n4898, B2 => n19244, C1 => n2418, C2 => 
                           n19238, A => n10045, ZN => n10042);
   U3289 : OAI221_X1 port map( B1 => n1840, B2 => n19196, C1 => n4219, C2 => 
                           n19190, A => n10047, ZN => n10040);
   U3290 : NOR4_X1 port map( A1 => n10013, A2 => n10014, A3 => n10015, A4 => 
                           n10016, ZN => n10012);
   U3291 : OAI221_X1 port map( B1 => n1840, B2 => n19395, C1 => n4219, C2 => 
                           n19389, A => n10025, ZN => n10013);
   U3292 : OAI221_X1 port map( B1 => n1914, B2 => n19467, C1 => n19463, C2 => 
                           n2215, A => n10017, ZN => n10016);
   U3293 : OAI221_X1 port map( B1 => n3343, B2 => n19419, C1 => n4827, C2 => 
                           n19413, A => n10022, ZN => n10014);
   U3294 : NOR4_X1 port map( A1 => n9973, A2 => n9974, A3 => n9975, A4 => n9976
                           , ZN => n9972);
   U3295 : OAI221_X1 port map( B1 => n1913, B2 => n19269, C1 => n19264, C2 => 
                           n2217, A => n9977, ZN => n9976);
   U3296 : OAI221_X1 port map( B1 => n4897, B2 => n19245, C1 => n2417, C2 => 
                           n19239, A => n9978, ZN => n9975);
   U3297 : OAI221_X1 port map( B1 => n1839, B2 => n19197, C1 => n4218, C2 => 
                           n19191, A => n9980, ZN => n9973);
   U3298 : NOR4_X1 port map( A1 => n9945, A2 => n9946, A3 => n9947, A4 => n9948
                           , ZN => n9944);
   U3299 : OAI221_X1 port map( B1 => n1839, B2 => n19396, C1 => n4218, C2 => 
                           n19390, A => n9958, ZN => n9945);
   U3300 : OAI221_X1 port map( B1 => n1913, B2 => n19468, C1 => n19463, C2 => 
                           n2218, A => n9949, ZN => n9948);
   U3301 : OAI221_X1 port map( B1 => n3342, B2 => n19420, C1 => n4826, C2 => 
                           n19414, A => n9955, ZN => n9946);
   U3302 : NOR4_X1 port map( A1 => n9906, A2 => n9907, A3 => n9908, A4 => n9909
                           , ZN => n9905);
   U3303 : OAI221_X1 port map( B1 => n1912, B2 => n19269, C1 => n19264, C2 => 
                           n2220, A => n9910, ZN => n9909);
   U3304 : OAI221_X1 port map( B1 => n4896, B2 => n19245, C1 => n2416, C2 => 
                           n19239, A => n9911, ZN => n9908);
   U3305 : OAI221_X1 port map( B1 => n1838, B2 => n19197, C1 => n4217, C2 => 
                           n19191, A => n9913, ZN => n9906);
   U3306 : NOR4_X1 port map( A1 => n9878, A2 => n9879, A3 => n9880, A4 => n9881
                           , ZN => n9877);
   U3307 : OAI221_X1 port map( B1 => n1838, B2 => n19396, C1 => n4217, C2 => 
                           n19390, A => n9890, ZN => n9878);
   U3308 : OAI221_X1 port map( B1 => n1912, B2 => n19468, C1 => n19463, C2 => 
                           n2221, A => n9882, ZN => n9881);
   U3309 : OAI221_X1 port map( B1 => n3341, B2 => n19420, C1 => n4825, C2 => 
                           n19414, A => n9887, ZN => n9879);
   U3310 : NOR4_X1 port map( A1 => n9838, A2 => n9839, A3 => n9840, A4 => n9841
                           , ZN => n9837);
   U3311 : OAI221_X1 port map( B1 => n1911, B2 => n19269, C1 => n19264, C2 => 
                           n2223, A => n9842, ZN => n9841);
   U3312 : OAI221_X1 port map( B1 => n4895, B2 => n19245, C1 => n2415, C2 => 
                           n19239, A => n9843, ZN => n9840);
   U3313 : OAI221_X1 port map( B1 => n1837, B2 => n19197, C1 => n4216, C2 => 
                           n19191, A => n9845, ZN => n9838);
   U3314 : NOR4_X1 port map( A1 => n9811, A2 => n9812, A3 => n9813, A4 => n9814
                           , ZN => n9810);
   U3315 : OAI221_X1 port map( B1 => n1837, B2 => n19396, C1 => n4216, C2 => 
                           n19390, A => n9823, ZN => n9811);
   U3316 : OAI221_X1 port map( B1 => n1911, B2 => n19468, C1 => n19463, C2 => 
                           n2224, A => n9815, ZN => n9814);
   U3317 : OAI221_X1 port map( B1 => n3340, B2 => n19420, C1 => n4824, C2 => 
                           n19414, A => n9820, ZN => n9812);
   U3318 : NOR4_X1 port map( A1 => n9771, A2 => n9772, A3 => n9773, A4 => n9774
                           , ZN => n9770);
   U3319 : OAI221_X1 port map( B1 => n1910, B2 => n19269, C1 => n19264, C2 => 
                           n2226, A => n9775, ZN => n9774);
   U3320 : OAI221_X1 port map( B1 => n4894, B2 => n19245, C1 => n2414, C2 => 
                           n19239, A => n9776, ZN => n9773);
   U3321 : OAI221_X1 port map( B1 => n1836, B2 => n19197, C1 => n4215, C2 => 
                           n19191, A => n9778, ZN => n9771);
   U3322 : NOR4_X1 port map( A1 => n9744, A2 => n9745, A3 => n9746, A4 => n9747
                           , ZN => n9743);
   U3323 : OAI221_X1 port map( B1 => n1836, B2 => n19396, C1 => n4215, C2 => 
                           n19390, A => n9756, ZN => n9744);
   U3324 : OAI221_X1 port map( B1 => n1910, B2 => n19468, C1 => n19463, C2 => 
                           n2227, A => n9748, ZN => n9747);
   U3325 : OAI221_X1 port map( B1 => n3339, B2 => n19420, C1 => n4823, C2 => 
                           n19414, A => n9753, ZN => n9745);
   U3326 : NOR4_X1 port map( A1 => n9704, A2 => n9705, A3 => n9706, A4 => n9707
                           , ZN => n9703);
   U3327 : OAI221_X1 port map( B1 => n1909, B2 => n19269, C1 => n19263, C2 => 
                           n2229, A => n9708, ZN => n9707);
   U3328 : OAI221_X1 port map( B1 => n4893, B2 => n19245, C1 => n2413, C2 => 
                           n19239, A => n9709, ZN => n9706);
   U3329 : OAI221_X1 port map( B1 => n1835, B2 => n19197, C1 => n4214, C2 => 
                           n19191, A => n9711, ZN => n9704);
   U3330 : NOR4_X1 port map( A1 => n9676, A2 => n9677, A3 => n9678, A4 => n9679
                           , ZN => n9675);
   U3331 : OAI221_X1 port map( B1 => n1835, B2 => n19396, C1 => n4214, C2 => 
                           n19390, A => n9688, ZN => n9676);
   U3332 : OAI221_X1 port map( B1 => n1909, B2 => n19468, C1 => n19462, C2 => 
                           n2230, A => n9680, ZN => n9679);
   U3333 : OAI221_X1 port map( B1 => n3338, B2 => n19420, C1 => n4822, C2 => 
                           n19414, A => n9685, ZN => n9677);
   U3334 : NOR4_X1 port map( A1 => n9637, A2 => n9638, A3 => n9639, A4 => n9640
                           , ZN => n9635);
   U3335 : OAI221_X1 port map( B1 => n1908, B2 => n19269, C1 => n19263, C2 => 
                           n2232, A => n9641, ZN => n9640);
   U3336 : OAI221_X1 port map( B1 => n4892, B2 => n19245, C1 => n2412, C2 => 
                           n19239, A => n9642, ZN => n9639);
   U3337 : OAI221_X1 port map( B1 => n1834, B2 => n19197, C1 => n4213, C2 => 
                           n19191, A => n9644, ZN => n9637);
   U3338 : NOR4_X1 port map( A1 => n9609, A2 => n9610, A3 => n9611, A4 => n9612
                           , ZN => n9608);
   U3339 : OAI221_X1 port map( B1 => n1834, B2 => n19396, C1 => n4213, C2 => 
                           n19390, A => n9621, ZN => n9609);
   U3340 : OAI221_X1 port map( B1 => n1908, B2 => n19468, C1 => n19462, C2 => 
                           n2233, A => n9613, ZN => n9612);
   U3341 : OAI221_X1 port map( B1 => n3337, B2 => n19420, C1 => n4821, C2 => 
                           n19414, A => n9618, ZN => n9610);
   U3342 : NOR4_X1 port map( A1 => n9569, A2 => n9570, A3 => n9571, A4 => n9572
                           , ZN => n9568);
   U3343 : OAI221_X1 port map( B1 => n1907, B2 => n19269, C1 => n19263, C2 => 
                           n2235, A => n9573, ZN => n9572);
   U3344 : OAI221_X1 port map( B1 => n4891, B2 => n19245, C1 => n2411, C2 => 
                           n19239, A => n9574, ZN => n9571);
   U3345 : OAI221_X1 port map( B1 => n1833, B2 => n19197, C1 => n4212, C2 => 
                           n19191, A => n9576, ZN => n9569);
   U3346 : NOR4_X1 port map( A1 => n9542, A2 => n9543, A3 => n9544, A4 => n9545
                           , ZN => n9541);
   U3347 : OAI221_X1 port map( B1 => n1833, B2 => n19396, C1 => n4212, C2 => 
                           n19390, A => n9554, ZN => n9542);
   U3348 : OAI221_X1 port map( B1 => n1907, B2 => n19468, C1 => n19462, C2 => 
                           n2236, A => n9546, ZN => n9545);
   U3349 : OAI221_X1 port map( B1 => n3336, B2 => n19420, C1 => n4820, C2 => 
                           n19414, A => n9551, ZN => n9543);
   U3350 : NOR4_X1 port map( A1 => n9502, A2 => n9503, A3 => n9504, A4 => n9505
                           , ZN => n9501);
   U3351 : OAI221_X1 port map( B1 => n1906, B2 => n19269, C1 => n19263, C2 => 
                           n2238, A => n9506, ZN => n9505);
   U3352 : OAI221_X1 port map( B1 => n4890, B2 => n19245, C1 => n2410, C2 => 
                           n19239, A => n9507, ZN => n9504);
   U3353 : OAI221_X1 port map( B1 => n1832, B2 => n19197, C1 => n4211, C2 => 
                           n19191, A => n9509, ZN => n9502);
   U3354 : NOR4_X1 port map( A1 => n9474, A2 => n9475, A3 => n9476, A4 => n9478
                           , ZN => n9473);
   U3355 : OAI221_X1 port map( B1 => n1832, B2 => n19396, C1 => n4211, C2 => 
                           n19390, A => n9487, ZN => n9474);
   U3356 : OAI221_X1 port map( B1 => n1906, B2 => n19468, C1 => n19462, C2 => 
                           n2239, A => n9479, ZN => n9478);
   U3357 : OAI221_X1 port map( B1 => n3335, B2 => n19420, C1 => n4819, C2 => 
                           n19414, A => n9484, ZN => n9475);
   U3358 : NOR4_X1 port map( A1 => n9435, A2 => n9436, A3 => n9437, A4 => n9438
                           , ZN => n9434);
   U3359 : OAI221_X1 port map( B1 => n1905, B2 => n19269, C1 => n19263, C2 => 
                           n2241, A => n9439, ZN => n9438);
   U3360 : OAI221_X1 port map( B1 => n4889, B2 => n19245, C1 => n2409, C2 => 
                           n19239, A => n9440, ZN => n9437);
   U3361 : OAI221_X1 port map( B1 => n1831, B2 => n19197, C1 => n4210, C2 => 
                           n19191, A => n9442, ZN => n9435);
   U3362 : NOR4_X1 port map( A1 => n9407, A2 => n9408, A3 => n9409, A4 => n9410
                           , ZN => n9406);
   U3363 : OAI221_X1 port map( B1 => n1831, B2 => n19396, C1 => n4210, C2 => 
                           n19390, A => n9419, ZN => n9407);
   U3364 : OAI221_X1 port map( B1 => n1905, B2 => n19468, C1 => n19462, C2 => 
                           n2242, A => n9411, ZN => n9410);
   U3365 : OAI221_X1 port map( B1 => n3334, B2 => n19420, C1 => n4818, C2 => 
                           n19414, A => n9416, ZN => n9408);
   U3366 : NOR4_X1 port map( A1 => n9367, A2 => n9368, A3 => n9369, A4 => n9370
                           , ZN => n9366);
   U3367 : OAI221_X1 port map( B1 => n1904, B2 => n19269, C1 => n19263, C2 => 
                           n2244, A => n9372, ZN => n9370);
   U3368 : OAI221_X1 port map( B1 => n4888, B2 => n19245, C1 => n2408, C2 => 
                           n19239, A => n9373, ZN => n9369);
   U3369 : OAI221_X1 port map( B1 => n1830, B2 => n19197, C1 => n4209, C2 => 
                           n19191, A => n9375, ZN => n9367);
   U3370 : NOR4_X1 port map( A1 => n9340, A2 => n9341, A3 => n9342, A4 => n9343
                           , ZN => n9339);
   U3371 : OAI221_X1 port map( B1 => n1830, B2 => n19396, C1 => n4209, C2 => 
                           n19390, A => n9352, ZN => n9340);
   U3372 : OAI221_X1 port map( B1 => n1904, B2 => n19468, C1 => n19462, C2 => 
                           n2245, A => n9344, ZN => n9343);
   U3373 : OAI221_X1 port map( B1 => n3333, B2 => n19420, C1 => n4817, C2 => 
                           n19414, A => n9349, ZN => n9341);
   U3374 : NOR4_X1 port map( A1 => n9300, A2 => n9301, A3 => n9302, A4 => n9303
                           , ZN => n9299);
   U3375 : OAI221_X1 port map( B1 => n1903, B2 => n19269, C1 => n19263, C2 => 
                           n2247, A => n9304, ZN => n9303);
   U3376 : OAI221_X1 port map( B1 => n4887, B2 => n19245, C1 => n2407, C2 => 
                           n19239, A => n9305, ZN => n9302);
   U3377 : OAI221_X1 port map( B1 => n1829, B2 => n19197, C1 => n4208, C2 => 
                           n19191, A => n9307, ZN => n9300);
   U3378 : NOR4_X1 port map( A1 => n9273, A2 => n9274, A3 => n9275, A4 => n9276
                           , ZN => n9272);
   U3379 : OAI221_X1 port map( B1 => n1829, B2 => n19396, C1 => n4208, C2 => 
                           n19390, A => n9285, ZN => n9273);
   U3380 : OAI221_X1 port map( B1 => n1903, B2 => n19468, C1 => n19462, C2 => 
                           n2248, A => n9277, ZN => n9276);
   U3381 : OAI221_X1 port map( B1 => n3332, B2 => n19420, C1 => n4816, C2 => 
                           n19414, A => n9282, ZN => n9274);
   U3382 : NOR4_X1 port map( A1 => n6993, A2 => n6994, A3 => n6995, A4 => n6996
                           , ZN => n6992);
   U3383 : OAI221_X1 port map( B1 => n1902, B2 => n19269, C1 => n19263, C2 => 
                           n2250, A => n6997, ZN => n6996);
   U3384 : OAI221_X1 port map( B1 => n4886, B2 => n19245, C1 => n2406, C2 => 
                           n19239, A => n6998, ZN => n6995);
   U3385 : OAI221_X1 port map( B1 => n1828, B2 => n19197, C1 => n4207, C2 => 
                           n19191, A => n7000, ZN => n6993);
   U3386 : NOR4_X1 port map( A1 => n6966, A2 => n6967, A3 => n6968, A4 => n6969
                           , ZN => n6965);
   U3387 : OAI221_X1 port map( B1 => n1828, B2 => n19396, C1 => n4207, C2 => 
                           n19390, A => n6978, ZN => n6966);
   U3388 : OAI221_X1 port map( B1 => n1902, B2 => n19468, C1 => n19462, C2 => 
                           n2251, A => n6970, ZN => n6969);
   U3389 : OAI221_X1 port map( B1 => n3331, B2 => n19420, C1 => n4815, C2 => 
                           n19414, A => n6975, ZN => n6967);
   U3390 : NOR4_X1 port map( A1 => n6926, A2 => n6927, A3 => n6928, A4 => n6929
                           , ZN => n6925);
   U3391 : OAI221_X1 port map( B1 => n1901, B2 => n19270, C1 => n19263, C2 => 
                           n2253, A => n6930, ZN => n6929);
   U3392 : OAI221_X1 port map( B1 => n4885, B2 => n19246, C1 => n2405, C2 => 
                           n19240, A => n6931, ZN => n6928);
   U3393 : OAI221_X1 port map( B1 => n1827, B2 => n19198, C1 => n4206, C2 => 
                           n19192, A => n6933, ZN => n6926);
   U3394 : NOR4_X1 port map( A1 => n6899, A2 => n6900, A3 => n6901, A4 => n6902
                           , ZN => n6898);
   U3395 : OAI221_X1 port map( B1 => n1827, B2 => n19397, C1 => n4206, C2 => 
                           n19391, A => n6911, ZN => n6899);
   U3396 : OAI221_X1 port map( B1 => n1901, B2 => n19469, C1 => n19462, C2 => 
                           n2254, A => n6903, ZN => n6902);
   U3397 : OAI221_X1 port map( B1 => n3330, B2 => n19421, C1 => n4814, C2 => 
                           n19415, A => n6908, ZN => n6900);
   U3398 : NOR4_X1 port map( A1 => n6859, A2 => n6860, A3 => n6861, A4 => n6862
                           , ZN => n6858);
   U3399 : OAI221_X1 port map( B1 => n1900, B2 => n19270, C1 => n19263, C2 => 
                           n2256, A => n6863, ZN => n6862);
   U3400 : OAI221_X1 port map( B1 => n4884, B2 => n19246, C1 => n2404, C2 => 
                           n19240, A => n6864, ZN => n6861);
   U3401 : OAI221_X1 port map( B1 => n1826, B2 => n19198, C1 => n4205, C2 => 
                           n19192, A => n6866, ZN => n6859);
   U3402 : NOR4_X1 port map( A1 => n6832, A2 => n6833, A3 => n6834, A4 => n6835
                           , ZN => n6831);
   U3403 : OAI221_X1 port map( B1 => n1826, B2 => n19397, C1 => n4205, C2 => 
                           n19391, A => n6844, ZN => n6832);
   U3404 : OAI221_X1 port map( B1 => n1900, B2 => n19469, C1 => n19462, C2 => 
                           n2257, A => n6836, ZN => n6835);
   U3405 : OAI221_X1 port map( B1 => n3329, B2 => n19421, C1 => n4813, C2 => 
                           n19415, A => n6841, ZN => n6833);
   U3406 : NOR4_X1 port map( A1 => n6792, A2 => n6793, A3 => n6794, A4 => n6795
                           , ZN => n6791);
   U3407 : OAI221_X1 port map( B1 => n1899, B2 => n19270, C1 => n19263, C2 => 
                           n2259, A => n6796, ZN => n6795);
   U3408 : OAI221_X1 port map( B1 => n4883, B2 => n19246, C1 => n2403, C2 => 
                           n19240, A => n6797, ZN => n6794);
   U3409 : OAI221_X1 port map( B1 => n1825, B2 => n19198, C1 => n4204, C2 => 
                           n19192, A => n6799, ZN => n6792);
   U3410 : NOR4_X1 port map( A1 => n6765, A2 => n6766, A3 => n6767, A4 => n6768
                           , ZN => n6764);
   U3411 : OAI221_X1 port map( B1 => n1825, B2 => n19397, C1 => n4204, C2 => 
                           n19391, A => n6777, ZN => n6765);
   U3412 : OAI221_X1 port map( B1 => n1899, B2 => n19469, C1 => n19462, C2 => 
                           n2260, A => n6769, ZN => n6768);
   U3413 : OAI221_X1 port map( B1 => n3328, B2 => n19421, C1 => n4812, C2 => 
                           n19415, A => n6774, ZN => n6766);
   U3414 : NOR4_X1 port map( A1 => n6725, A2 => n6726, A3 => n6727, A4 => n6728
                           , ZN => n6724);
   U3415 : OAI221_X1 port map( B1 => n1898, B2 => n19270, C1 => n19263, C2 => 
                           n2262, A => n6729, ZN => n6728);
   U3416 : OAI221_X1 port map( B1 => n4882, B2 => n19246, C1 => n2402, C2 => 
                           n19240, A => n6730, ZN => n6727);
   U3417 : OAI221_X1 port map( B1 => n1824, B2 => n19198, C1 => n4203, C2 => 
                           n19192, A => n6732, ZN => n6725);
   U3418 : NOR4_X1 port map( A1 => n6698, A2 => n6699, A3 => n6700, A4 => n6701
                           , ZN => n6697);
   U3419 : OAI221_X1 port map( B1 => n1824, B2 => n19397, C1 => n4203, C2 => 
                           n19391, A => n6710, ZN => n6698);
   U3420 : OAI221_X1 port map( B1 => n1898, B2 => n19469, C1 => n19462, C2 => 
                           n2263, A => n6702, ZN => n6701);
   U3421 : OAI221_X1 port map( B1 => n3327, B2 => n19421, C1 => n4811, C2 => 
                           n19415, A => n6707, ZN => n6699);
   U3422 : NOR4_X1 port map( A1 => n6658, A2 => n6659, A3 => n6660, A4 => n6661
                           , ZN => n6657);
   U3423 : OAI221_X1 port map( B1 => n1897, B2 => n19270, C1 => n19262, C2 => 
                           n2265, A => n6662, ZN => n6661);
   U3424 : OAI221_X1 port map( B1 => n4881, B2 => n19246, C1 => n2401, C2 => 
                           n19240, A => n6663, ZN => n6660);
   U3425 : OAI221_X1 port map( B1 => n1823, B2 => n19198, C1 => n4202, C2 => 
                           n19192, A => n6665, ZN => n6658);
   U3426 : NOR4_X1 port map( A1 => n6630, A2 => n6631, A3 => n6632, A4 => n6633
                           , ZN => n6629);
   U3427 : OAI221_X1 port map( B1 => n1823, B2 => n19397, C1 => n4202, C2 => 
                           n19391, A => n6642, ZN => n6630);
   U3428 : OAI221_X1 port map( B1 => n1897, B2 => n19469, C1 => n19461, C2 => 
                           n2266, A => n6634, ZN => n6633);
   U3429 : OAI221_X1 port map( B1 => n3326, B2 => n19421, C1 => n4810, C2 => 
                           n19415, A => n6639, ZN => n6631);
   U3430 : NOR4_X1 port map( A1 => n6591, A2 => n6592, A3 => n6593, A4 => n6594
                           , ZN => n6590);
   U3431 : OAI221_X1 port map( B1 => n1896, B2 => n19270, C1 => n19262, C2 => 
                           n2268, A => n6595, ZN => n6594);
   U3432 : OAI221_X1 port map( B1 => n4880, B2 => n19246, C1 => n2400, C2 => 
                           n19240, A => n6596, ZN => n6593);
   U3433 : OAI221_X1 port map( B1 => n1822, B2 => n19198, C1 => n4201, C2 => 
                           n19192, A => n6598, ZN => n6591);
   U3434 : NOR4_X1 port map( A1 => n6564, A2 => n6565, A3 => n6566, A4 => n6567
                           , ZN => n6563);
   U3435 : OAI221_X1 port map( B1 => n1822, B2 => n19397, C1 => n4201, C2 => 
                           n19391, A => n6576, ZN => n6564);
   U3436 : OAI221_X1 port map( B1 => n1896, B2 => n19469, C1 => n19461, C2 => 
                           n2269, A => n6568, ZN => n6567);
   U3437 : OAI221_X1 port map( B1 => n3325, B2 => n19421, C1 => n4809, C2 => 
                           n19415, A => n6573, ZN => n6565);
   U3438 : NOR4_X1 port map( A1 => n6525, A2 => n6526, A3 => n6527, A4 => n6528
                           , ZN => n6524);
   U3439 : OAI221_X1 port map( B1 => n1895, B2 => n19270, C1 => n19262, C2 => 
                           n2271, A => n6529, ZN => n6528);
   U3440 : OAI221_X1 port map( B1 => n4879, B2 => n19246, C1 => n2399, C2 => 
                           n19240, A => n6530, ZN => n6527);
   U3441 : OAI221_X1 port map( B1 => n1821, B2 => n19198, C1 => n4200, C2 => 
                           n19192, A => n6532, ZN => n6525);
   U3442 : NOR4_X1 port map( A1 => n6498, A2 => n6499, A3 => n6500, A4 => n6501
                           , ZN => n6497);
   U3443 : OAI221_X1 port map( B1 => n1821, B2 => n19397, C1 => n4200, C2 => 
                           n19391, A => n6510, ZN => n6498);
   U3444 : OAI221_X1 port map( B1 => n1895, B2 => n19469, C1 => n19461, C2 => 
                           n2272, A => n6502, ZN => n6501);
   U3445 : OAI221_X1 port map( B1 => n3324, B2 => n19421, C1 => n4808, C2 => 
                           n19415, A => n6507, ZN => n6499);
   U3446 : NOR4_X1 port map( A1 => n6459, A2 => n6460, A3 => n6461, A4 => n6462
                           , ZN => n6458);
   U3447 : OAI221_X1 port map( B1 => n1894, B2 => n19270, C1 => n19262, C2 => 
                           n2274, A => n6463, ZN => n6462);
   U3448 : OAI221_X1 port map( B1 => n4878, B2 => n19246, C1 => n2398, C2 => 
                           n19240, A => n6464, ZN => n6461);
   U3449 : OAI221_X1 port map( B1 => n1820, B2 => n19198, C1 => n4199, C2 => 
                           n19192, A => n6466, ZN => n6459);
   U3450 : NOR4_X1 port map( A1 => n6432, A2 => n6433, A3 => n6434, A4 => n6435
                           , ZN => n6431);
   U3451 : OAI221_X1 port map( B1 => n1820, B2 => n19397, C1 => n4199, C2 => 
                           n19391, A => n6444, ZN => n6432);
   U3452 : OAI221_X1 port map( B1 => n1894, B2 => n19469, C1 => n19461, C2 => 
                           n2275, A => n6436, ZN => n6435);
   U3453 : OAI221_X1 port map( B1 => n3323, B2 => n19421, C1 => n4807, C2 => 
                           n19415, A => n6441, ZN => n6433);
   U3454 : NOR4_X1 port map( A1 => n6393, A2 => n6394, A3 => n6395, A4 => n6396
                           , ZN => n6392);
   U3455 : OAI221_X1 port map( B1 => n1893, B2 => n19270, C1 => n19262, C2 => 
                           n2277, A => n6397, ZN => n6396);
   U3456 : OAI221_X1 port map( B1 => n4877, B2 => n19246, C1 => n2397, C2 => 
                           n19240, A => n6398, ZN => n6395);
   U3457 : OAI221_X1 port map( B1 => n1819, B2 => n19198, C1 => n4198, C2 => 
                           n19192, A => n6400, ZN => n6393);
   U3458 : NOR4_X1 port map( A1 => n6366, A2 => n6367, A3 => n6368, A4 => n6369
                           , ZN => n6365);
   U3459 : OAI221_X1 port map( B1 => n1819, B2 => n19397, C1 => n4198, C2 => 
                           n19391, A => n6378, ZN => n6366);
   U3460 : OAI221_X1 port map( B1 => n1893, B2 => n19469, C1 => n19461, C2 => 
                           n2278, A => n6370, ZN => n6369);
   U3461 : OAI221_X1 port map( B1 => n3322, B2 => n19421, C1 => n4806, C2 => 
                           n19415, A => n6375, ZN => n6367);
   U3462 : NOR4_X1 port map( A1 => n6327, A2 => n6328, A3 => n6329, A4 => n6330
                           , ZN => n6326);
   U3463 : OAI221_X1 port map( B1 => n1892, B2 => n19270, C1 => n19262, C2 => 
                           n2280, A => n6331, ZN => n6330);
   U3464 : OAI221_X1 port map( B1 => n4876, B2 => n19246, C1 => n2396, C2 => 
                           n19240, A => n6332, ZN => n6329);
   U3465 : OAI221_X1 port map( B1 => n1818, B2 => n19198, C1 => n4197, C2 => 
                           n19192, A => n6334, ZN => n6327);
   U3466 : NOR4_X1 port map( A1 => n6300, A2 => n6301, A3 => n6302, A4 => n6303
                           , ZN => n6299);
   U3467 : OAI221_X1 port map( B1 => n1818, B2 => n19397, C1 => n4197, C2 => 
                           n19391, A => n6312, ZN => n6300);
   U3468 : OAI221_X1 port map( B1 => n1892, B2 => n19469, C1 => n19461, C2 => 
                           n2281, A => n6304, ZN => n6303);
   U3469 : OAI221_X1 port map( B1 => n3321, B2 => n19421, C1 => n4805, C2 => 
                           n19415, A => n6309, ZN => n6301);
   U3470 : NOR4_X1 port map( A1 => n6261, A2 => n6262, A3 => n6263, A4 => n6264
                           , ZN => n6260);
   U3471 : OAI221_X1 port map( B1 => n1891, B2 => n19270, C1 => n19262, C2 => 
                           n2283, A => n6265, ZN => n6264);
   U3472 : OAI221_X1 port map( B1 => n4875, B2 => n19246, C1 => n2395, C2 => 
                           n19240, A => n6266, ZN => n6263);
   U3473 : OAI221_X1 port map( B1 => n1817, B2 => n19198, C1 => n4196, C2 => 
                           n19192, A => n6268, ZN => n6261);
   U3474 : NOR4_X1 port map( A1 => n6234, A2 => n6235, A3 => n6236, A4 => n6237
                           , ZN => n6233);
   U3475 : OAI221_X1 port map( B1 => n1817, B2 => n19397, C1 => n4196, C2 => 
                           n19391, A => n6246, ZN => n6234);
   U3476 : OAI221_X1 port map( B1 => n1891, B2 => n19469, C1 => n19461, C2 => 
                           n2284, A => n6238, ZN => n6237);
   U3477 : OAI221_X1 port map( B1 => n3320, B2 => n19421, C1 => n4804, C2 => 
                           n19415, A => n6243, ZN => n6235);
   U3478 : NOR4_X1 port map( A1 => n6195, A2 => n6196, A3 => n6197, A4 => n6198
                           , ZN => n6194);
   U3479 : OAI221_X1 port map( B1 => n1890, B2 => n19270, C1 => n19262, C2 => 
                           n2286, A => n6199, ZN => n6198);
   U3480 : OAI221_X1 port map( B1 => n4874, B2 => n19246, C1 => n2394, C2 => 
                           n19240, A => n6200, ZN => n6197);
   U3481 : OAI221_X1 port map( B1 => n1816, B2 => n19198, C1 => n4195, C2 => 
                           n19192, A => n6202, ZN => n6195);
   U3482 : NOR4_X1 port map( A1 => n6168, A2 => n6169, A3 => n6170, A4 => n6171
                           , ZN => n6167);
   U3483 : OAI221_X1 port map( B1 => n1816, B2 => n19397, C1 => n4195, C2 => 
                           n19391, A => n6180, ZN => n6168);
   U3484 : OAI221_X1 port map( B1 => n1890, B2 => n19469, C1 => n19461, C2 => 
                           n2287, A => n6172, ZN => n6171);
   U3485 : OAI221_X1 port map( B1 => n3319, B2 => n19421, C1 => n4803, C2 => 
                           n19415, A => n6177, ZN => n6169);
   U3486 : NOR4_X1 port map( A1 => n6129, A2 => n6130, A3 => n6131, A4 => n6132
                           , ZN => n6128);
   U3487 : OAI221_X1 port map( B1 => n1889, B2 => n19271, C1 => n19262, C2 => 
                           n2289, A => n6133, ZN => n6132);
   U3488 : OAI221_X1 port map( B1 => n4873, B2 => n19247, C1 => n2393, C2 => 
                           n19241, A => n6134, ZN => n6131);
   U3489 : OAI221_X1 port map( B1 => n1815, B2 => n19199, C1 => n4194, C2 => 
                           n19193, A => n6136, ZN => n6129);
   U3490 : NOR4_X1 port map( A1 => n6102, A2 => n6103, A3 => n6104, A4 => n6105
                           , ZN => n6101);
   U3491 : OAI221_X1 port map( B1 => n1815, B2 => n19398, C1 => n4194, C2 => 
                           n19392, A => n6114, ZN => n6102);
   U3492 : OAI221_X1 port map( B1 => n1889, B2 => n19470, C1 => n19461, C2 => 
                           n2290, A => n6106, ZN => n6105);
   U3493 : OAI221_X1 port map( B1 => n3318, B2 => n19422, C1 => n4802, C2 => 
                           n19416, A => n6111, ZN => n6103);
   U3494 : NOR4_X1 port map( A1 => n6063, A2 => n6064, A3 => n6065, A4 => n6066
                           , ZN => n6062);
   U3495 : OAI221_X1 port map( B1 => n1888, B2 => n19271, C1 => n19262, C2 => 
                           n2292, A => n6067, ZN => n6066);
   U3496 : OAI221_X1 port map( B1 => n4872, B2 => n19247, C1 => n2392, C2 => 
                           n19241, A => n6068, ZN => n6065);
   U3497 : OAI221_X1 port map( B1 => n1814, B2 => n19199, C1 => n4193, C2 => 
                           n19193, A => n6070, ZN => n6063);
   U3498 : NOR4_X1 port map( A1 => n6036, A2 => n6037, A3 => n6038, A4 => n6039
                           , ZN => n6034);
   U3499 : OAI221_X1 port map( B1 => n1814, B2 => n19398, C1 => n4193, C2 => 
                           n19392, A => n6048, ZN => n6036);
   U3500 : OAI221_X1 port map( B1 => n1888, B2 => n19470, C1 => n19461, C2 => 
                           n2293, A => n6040, ZN => n6039);
   U3501 : OAI221_X1 port map( B1 => n3317, B2 => n19422, C1 => n4801, C2 => 
                           n19416, A => n6045, ZN => n6037);
   U3502 : NOR4_X1 port map( A1 => n5995, A2 => n5996, A3 => n5997, A4 => n5998
                           , ZN => n5994);
   U3503 : OAI221_X1 port map( B1 => n1887, B2 => n19271, C1 => n19262, C2 => 
                           n2295, A => n5999, ZN => n5998);
   U3504 : OAI221_X1 port map( B1 => n4871, B2 => n19247, C1 => n2391, C2 => 
                           n19241, A => n6000, ZN => n5997);
   U3505 : OAI221_X1 port map( B1 => n1813, B2 => n19199, C1 => n4192, C2 => 
                           n19193, A => n6002, ZN => n5995);
   U3506 : NOR4_X1 port map( A1 => n5967, A2 => n5969, A3 => n5970, A4 => n5971
                           , ZN => n5965);
   U3507 : OAI221_X1 port map( B1 => n1813, B2 => n19398, C1 => n4192, C2 => 
                           n19392, A => n5980, ZN => n5967);
   U3508 : OAI221_X1 port map( B1 => n1887, B2 => n19470, C1 => n19461, C2 => 
                           n2296, A => n5972, ZN => n5971);
   U3509 : OAI221_X1 port map( B1 => n3316, B2 => n19422, C1 => n4800, C2 => 
                           n19416, A => n5977, ZN => n5969);
   U3510 : NOR4_X1 port map( A1 => n5927, A2 => n5928, A3 => n5929, A4 => n5930
                           , ZN => n5926);
   U3511 : OAI221_X1 port map( B1 => n1886, B2 => n19271, C1 => n19262, C2 => 
                           n2298, A => n5931, ZN => n5930);
   U3512 : OAI221_X1 port map( B1 => n4870, B2 => n19247, C1 => n2390, C2 => 
                           n19241, A => n5932, ZN => n5929);
   U3513 : OAI221_X1 port map( B1 => n1812, B2 => n19199, C1 => n4191, C2 => 
                           n19193, A => n5934, ZN => n5927);
   U3514 : NOR4_X1 port map( A1 => n5899, A2 => n5900, A3 => n5902, A4 => n5903
                           , ZN => n5898);
   U3515 : OAI221_X1 port map( B1 => n1812, B2 => n19398, C1 => n4191, C2 => 
                           n19392, A => n5912, ZN => n5899);
   U3516 : OAI221_X1 port map( B1 => n1886, B2 => n19470, C1 => n19461, C2 => 
                           n2299, A => n5904, ZN => n5903);
   U3517 : OAI221_X1 port map( B1 => n3315, B2 => n19422, C1 => n4799, C2 => 
                           n19416, A => n5909, ZN => n5900);
   U3518 : NOR4_X1 port map( A1 => n5860, A2 => n5861, A3 => n5862, A4 => n5863
                           , ZN => n5859);
   U3519 : OAI221_X1 port map( B1 => n1885, B2 => n19271, C1 => n19261, C2 => 
                           n2301, A => n5864, ZN => n5863);
   U3520 : OAI221_X1 port map( B1 => n4869, B2 => n19247, C1 => n2389, C2 => 
                           n19241, A => n5865, ZN => n5862);
   U3521 : OAI221_X1 port map( B1 => n1811, B2 => n19199, C1 => n4190, C2 => 
                           n19193, A => n5867, ZN => n5860);
   U3522 : NOR4_X1 port map( A1 => n5832, A2 => n5833, A3 => n5834, A4 => n5836
                           , ZN => n5831);
   U3523 : OAI221_X1 port map( B1 => n1811, B2 => n19398, C1 => n4190, C2 => 
                           n19392, A => n5845, ZN => n5832);
   U3524 : OAI221_X1 port map( B1 => n1885, B2 => n19470, C1 => n19460, C2 => 
                           n2302, A => n5837, ZN => n5836);
   U3525 : OAI221_X1 port map( B1 => n3314, B2 => n19422, C1 => n4798, C2 => 
                           n19416, A => n5842, ZN => n5833);
   U3526 : NOR4_X1 port map( A1 => n5793, A2 => n5794, A3 => n5795, A4 => n5796
                           , ZN => n5792);
   U3527 : OAI221_X1 port map( B1 => n1884, B2 => n19271, C1 => n19261, C2 => 
                           n2304, A => n5797, ZN => n5796);
   U3528 : OAI221_X1 port map( B1 => n4868, B2 => n19247, C1 => n2388, C2 => 
                           n19241, A => n5798, ZN => n5795);
   U3529 : OAI221_X1 port map( B1 => n1810, B2 => n19199, C1 => n4189, C2 => 
                           n19193, A => n5800, ZN => n5793);
   U3530 : NOR4_X1 port map( A1 => n5760, A2 => n5761, A3 => n5762, A4 => n5768
                           , ZN => n5759);
   U3531 : OAI221_X1 port map( B1 => n1810, B2 => n19398, C1 => n4189, C2 => 
                           n19392, A => n5778, ZN => n5760);
   U3532 : OAI221_X1 port map( B1 => n1884, B2 => n19470, C1 => n19460, C2 => 
                           n2305, A => n5770, ZN => n5768);
   U3533 : OAI221_X1 port map( B1 => n3313, B2 => n19422, C1 => n4797, C2 => 
                           n19416, A => n5775, ZN => n5761);
   U3534 : NOR4_X1 port map( A1 => n5721, A2 => n5722, A3 => n5723, A4 => n5724
                           , ZN => n5720);
   U3535 : OAI221_X1 port map( B1 => n1883, B2 => n19271, C1 => n19261, C2 => 
                           n2307, A => n5725, ZN => n5724);
   U3536 : OAI221_X1 port map( B1 => n4867, B2 => n19247, C1 => n2387, C2 => 
                           n19241, A => n5726, ZN => n5723);
   U3537 : OAI221_X1 port map( B1 => n1809, B2 => n19199, C1 => n4188, C2 => 
                           n19193, A => n5728, ZN => n5721);
   U3538 : NOR4_X1 port map( A1 => n5690, A2 => n5691, A3 => n5692, A4 => n5693
                           , ZN => n5689);
   U3539 : OAI221_X1 port map( B1 => n1809, B2 => n19398, C1 => n4188, C2 => 
                           n19392, A => n5706, ZN => n5690);
   U3540 : OAI221_X1 port map( B1 => n1883, B2 => n19470, C1 => n19460, C2 => 
                           n2308, A => n5697, ZN => n5693);
   U3541 : OAI221_X1 port map( B1 => n3312, B2 => n19422, C1 => n4796, C2 => 
                           n19416, A => n5703, ZN => n5691);
   U3542 : NOR4_X1 port map( A1 => n5651, A2 => n5652, A3 => n5653, A4 => n5654
                           , ZN => n5650);
   U3543 : OAI221_X1 port map( B1 => n1882, B2 => n19271, C1 => n19261, C2 => 
                           n2310, A => n5655, ZN => n5654);
   U3544 : OAI221_X1 port map( B1 => n4866, B2 => n19247, C1 => n2386, C2 => 
                           n19241, A => n5656, ZN => n5653);
   U3545 : OAI221_X1 port map( B1 => n1808, B2 => n19199, C1 => n4187, C2 => 
                           n19193, A => n5658, ZN => n5651);
   U3546 : NOR4_X1 port map( A1 => n5622, A2 => n5623, A3 => n5624, A4 => n5625
                           , ZN => n5621);
   U3547 : OAI221_X1 port map( B1 => n1808, B2 => n19398, C1 => n4187, C2 => 
                           n19392, A => n5636, ZN => n5622);
   U3548 : OAI221_X1 port map( B1 => n1882, B2 => n19470, C1 => n19460, C2 => 
                           n2311, A => n5626, ZN => n5625);
   U3549 : OAI221_X1 port map( B1 => n3311, B2 => n19422, C1 => n4795, C2 => 
                           n19416, A => n5633, ZN => n5623);
   U3550 : NOR4_X1 port map( A1 => n5583, A2 => n5584, A3 => n5585, A4 => n5586
                           , ZN => n5582);
   U3551 : OAI221_X1 port map( B1 => n1881, B2 => n19271, C1 => n19261, C2 => 
                           n2313, A => n5587, ZN => n5586);
   U3552 : OAI221_X1 port map( B1 => n4865, B2 => n19247, C1 => n2385, C2 => 
                           n19241, A => n5588, ZN => n5585);
   U3553 : OAI221_X1 port map( B1 => n1807, B2 => n19199, C1 => n4186, C2 => 
                           n19193, A => n5590, ZN => n5583);
   U3554 : NOR4_X1 port map( A1 => n5553, A2 => n5554, A3 => n5555, A4 => n5556
                           , ZN => n5552);
   U3555 : OAI221_X1 port map( B1 => n1807, B2 => n19398, C1 => n4186, C2 => 
                           n19392, A => n5568, ZN => n5553);
   U3556 : OAI221_X1 port map( B1 => n1881, B2 => n19470, C1 => n19460, C2 => 
                           n2314, A => n5557, ZN => n5556);
   U3557 : OAI221_X1 port map( B1 => n3310, B2 => n19422, C1 => n4794, C2 => 
                           n19416, A => n5565, ZN => n5554);
   U3558 : NOR4_X1 port map( A1 => n5514, A2 => n5515, A3 => n5516, A4 => n5517
                           , ZN => n5513);
   U3559 : OAI221_X1 port map( B1 => n1880, B2 => n19271, C1 => n19261, C2 => 
                           n2316, A => n5518, ZN => n5517);
   U3560 : OAI221_X1 port map( B1 => n4864, B2 => n19247, C1 => n2384, C2 => 
                           n19241, A => n5519, ZN => n5516);
   U3561 : OAI221_X1 port map( B1 => n1806, B2 => n19199, C1 => n4185, C2 => 
                           n19193, A => n5521, ZN => n5514);
   U3562 : NOR4_X1 port map( A1 => n5484, A2 => n5485, A3 => n5486, A4 => n5487
                           , ZN => n5483);
   U3563 : OAI221_X1 port map( B1 => n1806, B2 => n19398, C1 => n4185, C2 => 
                           n19392, A => n5499, ZN => n5484);
   U3564 : OAI221_X1 port map( B1 => n1880, B2 => n19470, C1 => n19460, C2 => 
                           n2317, A => n5488, ZN => n5487);
   U3565 : OAI221_X1 port map( B1 => n3309, B2 => n19422, C1 => n4793, C2 => 
                           n19416, A => n5496, ZN => n5485);
   U3566 : NOR4_X1 port map( A1 => n5445, A2 => n5446, A3 => n5447, A4 => n5448
                           , ZN => n5444);
   U3567 : OAI221_X1 port map( B1 => n1879, B2 => n19271, C1 => n19261, C2 => 
                           n2319, A => n5449, ZN => n5448);
   U3568 : OAI221_X1 port map( B1 => n4863, B2 => n19247, C1 => n2383, C2 => 
                           n19241, A => n5450, ZN => n5447);
   U3569 : OAI221_X1 port map( B1 => n1805, B2 => n19199, C1 => n4184, C2 => 
                           n19193, A => n5452, ZN => n5445);
   U3570 : NOR4_X1 port map( A1 => n5416, A2 => n5417, A3 => n5418, A4 => n5419
                           , ZN => n5415);
   U3571 : OAI221_X1 port map( B1 => n1805, B2 => n19398, C1 => n4184, C2 => 
                           n19392, A => n5430, ZN => n5416);
   U3572 : OAI221_X1 port map( B1 => n1879, B2 => n19470, C1 => n19460, C2 => 
                           n2320, A => n5420, ZN => n5419);
   U3573 : OAI221_X1 port map( B1 => n3308, B2 => n19422, C1 => n4792, C2 => 
                           n19416, A => n5427, ZN => n5417);
   U3574 : NOR4_X1 port map( A1 => n5377, A2 => n5378, A3 => n5379, A4 => n5380
                           , ZN => n5376);
   U3575 : OAI221_X1 port map( B1 => n1878, B2 => n19271, C1 => n19261, C2 => 
                           n2322, A => n5381, ZN => n5380);
   U3576 : OAI221_X1 port map( B1 => n4862, B2 => n19247, C1 => n2382, C2 => 
                           n19241, A => n5382, ZN => n5379);
   U3577 : OAI221_X1 port map( B1 => n1804, B2 => n19199, C1 => n4183, C2 => 
                           n19193, A => n5384, ZN => n5377);
   U3578 : NOR4_X1 port map( A1 => n5346, A2 => n5347, A3 => n5348, A4 => n5349
                           , ZN => n5345);
   U3579 : OAI221_X1 port map( B1 => n1804, B2 => n19398, C1 => n4183, C2 => 
                           n19392, A => n5362, ZN => n5346);
   U3580 : OAI221_X1 port map( B1 => n1878, B2 => n19470, C1 => n19460, C2 => 
                           n2323, A => n5350, ZN => n5349);
   U3581 : OAI221_X1 port map( B1 => n3307, B2 => n19422, C1 => n4791, C2 => 
                           n19416, A => n5358, ZN => n5347);
   U3582 : NOR2_X1 port map( A1 => fill, A2 => spill, ZN => n2092);
   U3583 : OAI222_X1 port map( A1 => n1758, A2 => n19071, B1 => n3798, B2 => 
                           n19065, C1 => n3732, C2 => n19059, ZN => n6814);
   U3584 : OAI21_X1 port map( B1 => n11661, B2 => n11557, A => n20354, ZN => 
                           n3033);
   U3585 : INV_X1 port map( A => rd1, ZN => n11661);
   U3586 : AOI211_X1 port map( C1 => registers_4_38_port, C2 => n18981, A => 
                           n6819, B => n6820, ZN => n6809);
   U3587 : OAI221_X1 port map( B1 => n3599, B2 => n18963, C1 => n18957, C2 => 
                           n2725, A => n6821, ZN => n6819);
   U3588 : OAI22_X1 port map( A1 => n4949, A2 => n18975, B1 => n5015, B2 => 
                           n18969, ZN => n6820);
   U3589 : AOI22_X1 port map( A1 => n18951, A2 => n18116, B1 => n18945, B2 => 
                           n17696, ZN => n6821);
   U3590 : XNOR2_X1 port map( A => n11737, B => n11738, ZN => n1871);
   U3591 : XNOR2_X1 port map( A => count3(1), B => n11681, ZN => n11738);
   U3592 : OAI221_X1 port map( B1 => n1815, B2 => n19054, C1 => n5272, C2 => 
                           n19048, A => n6151, ZN => n6149);
   U3593 : AOI22_X1 port map( A1 => n19042, A2 => n17876, B1 => n19036, B2 => 
                           n17756, ZN => n6151);
   U3594 : OAI221_X1 port map( B1 => n1814, B2 => n19054, C1 => n5271, C2 => 
                           n19048, A => n6085, ZN => n6083);
   U3595 : AOI22_X1 port map( A1 => n19042, A2 => n17877, B1 => n19036, B2 => 
                           n17757, ZN => n6085);
   U3596 : OAI221_X1 port map( B1 => n1813, B2 => n19054, C1 => n5270, C2 => 
                           n19048, A => n6017, ZN => n6015);
   U3597 : AOI22_X1 port map( A1 => n19042, A2 => n17878, B1 => n19036, B2 => 
                           n17758, ZN => n6017);
   U3598 : OAI221_X1 port map( B1 => n1812, B2 => n19054, C1 => n5269, C2 => 
                           n19048, A => n5949, ZN => n5947);
   U3599 : AOI22_X1 port map( A1 => n19042, A2 => n17879, B1 => n19036, B2 => 
                           n17759, ZN => n5949);
   U3600 : OAI221_X1 port map( B1 => n1811, B2 => n19054, C1 => n5268, C2 => 
                           n19048, A => n5882, ZN => n5880);
   U3601 : AOI22_X1 port map( A1 => n19042, A2 => n17880, B1 => n19036, B2 => 
                           n17760, ZN => n5882);
   U3602 : OAI221_X1 port map( B1 => n1810, B2 => n19054, C1 => n5267, C2 => 
                           n19048, A => n5815, ZN => n5813);
   U3603 : AOI22_X1 port map( A1 => n19042, A2 => n17881, B1 => n19036, B2 => 
                           n17761, ZN => n5815);
   U3604 : OAI221_X1 port map( B1 => n1809, B2 => n19054, C1 => n5266, C2 => 
                           n19048, A => n5743, ZN => n5741);
   U3605 : AOI22_X1 port map( A1 => n19042, A2 => n17882, B1 => n19036, B2 => 
                           n17762, ZN => n5743);
   U3606 : OAI221_X1 port map( B1 => n1808, B2 => n19054, C1 => n5265, C2 => 
                           n19048, A => n5673, ZN => n5671);
   U3607 : AOI22_X1 port map( A1 => n19042, A2 => n17883, B1 => n19036, B2 => 
                           n17763, ZN => n5673);
   U3608 : OAI221_X1 port map( B1 => n1807, B2 => n19054, C1 => n5264, C2 => 
                           n19048, A => n5605, ZN => n5603);
   U3609 : AOI22_X1 port map( A1 => n19042, A2 => n17884, B1 => n19036, B2 => 
                           n17764, ZN => n5605);
   U3610 : OAI221_X1 port map( B1 => n1806, B2 => n19054, C1 => n5263, C2 => 
                           n19048, A => n5536, ZN => n5534);
   U3611 : AOI22_X1 port map( A1 => n19042, A2 => n17885, B1 => n19036, B2 => 
                           n17765, ZN => n5536);
   U3612 : OAI221_X1 port map( B1 => n1805, B2 => n19054, C1 => n5262, C2 => 
                           n19048, A => n5467, ZN => n5465);
   U3613 : AOI22_X1 port map( A1 => n19042, A2 => n17886, B1 => n19036, B2 => 
                           n17766, ZN => n5467);
   U3614 : OAI221_X1 port map( B1 => n1804, B2 => n19054, C1 => n5261, C2 => 
                           n19048, A => n5399, ZN => n5397);
   U3615 : AOI22_X1 port map( A1 => n19042, A2 => n17887, B1 => n19036, B2 => 
                           n17767, ZN => n5399);
   U3616 : OAI221_X1 port map( B1 => n1851, B2 => n19051, C1 => n5696, C2 => 
                           n19045, A => n10803, ZN => n10800);
   U3617 : AOI22_X1 port map( A1 => n19039, A2 => n17888, B1 => n19033, B2 => 
                           n17768, ZN => n10803);
   U3618 : OAI221_X1 port map( B1 => n1850, B2 => n19051, C1 => n5695, C2 => 
                           n19045, A => n10735, ZN => n10733);
   U3619 : AOI22_X1 port map( A1 => n19039, A2 => n17889, B1 => n19033, B2 => 
                           n17769, ZN => n10735);
   U3620 : OAI221_X1 port map( B1 => n1849, B2 => n19051, C1 => n5694, C2 => 
                           n19045, A => n10668, ZN => n10666);
   U3621 : AOI22_X1 port map( A1 => n19039, A2 => n17890, B1 => n19033, B2 => 
                           n17770, ZN => n10668);
   U3622 : OAI221_X1 port map( B1 => n1848, B2 => n19051, C1 => n5629, C2 => 
                           n19045, A => n10601, ZN => n10599);
   U3623 : AOI22_X1 port map( A1 => n19039, A2 => n17891, B1 => n19033, B2 => 
                           n17771, ZN => n10601);
   U3624 : OAI221_X1 port map( B1 => n1847, B2 => n19051, C1 => n5627, C2 => 
                           n19045, A => n10533, ZN => n10531);
   U3625 : AOI22_X1 port map( A1 => n19039, A2 => n17892, B1 => n19033, B2 => 
                           n17772, ZN => n10533);
   U3626 : OAI221_X1 port map( B1 => n1846, B2 => n19051, C1 => n5562, C2 => 
                           n19045, A => n10466, ZN => n10464);
   U3627 : AOI22_X1 port map( A1 => n19039, A2 => n17893, B1 => n19033, B2 => 
                           n17773, ZN => n10466);
   U3628 : OAI221_X1 port map( B1 => n1845, B2 => n19051, C1 => n5560, C2 => 
                           n19045, A => n10399, ZN => n10397);
   U3629 : AOI22_X1 port map( A1 => n19039, A2 => n17894, B1 => n19033, B2 => 
                           n17774, ZN => n10399);
   U3630 : OAI221_X1 port map( B1 => n1844, B2 => n19051, C1 => n5559, C2 => 
                           n19045, A => n10332, ZN => n10330);
   U3631 : AOI22_X1 port map( A1 => n19039, A2 => n17895, B1 => n19033, B2 => 
                           n17775, ZN => n10332);
   U3632 : OAI221_X1 port map( B1 => n1843, B2 => n19051, C1 => n5494, C2 => 
                           n19045, A => n10264, ZN => n10262);
   U3633 : AOI22_X1 port map( A1 => n19039, A2 => n17896, B1 => n19033, B2 => 
                           n17776, ZN => n10264);
   U3634 : OAI221_X1 port map( B1 => n1842, B2 => n19051, C1 => n5492, C2 => 
                           n19045, A => n10197, ZN => n10195);
   U3635 : AOI22_X1 port map( A1 => n19039, A2 => n17897, B1 => n19033, B2 => 
                           n17777, ZN => n10197);
   U3636 : OAI221_X1 port map( B1 => n1841, B2 => n19051, C1 => n5491, C2 => 
                           n19045, A => n10130, ZN => n10128);
   U3637 : AOI22_X1 port map( A1 => n19039, A2 => n17898, B1 => n19033, B2 => 
                           n17778, ZN => n10130);
   U3638 : OAI221_X1 port map( B1 => n1840, B2 => n19051, C1 => n5426, C2 => 
                           n19045, A => n10063, ZN => n10061);
   U3639 : AOI22_X1 port map( A1 => n19039, A2 => n17899, B1 => n19033, B2 => 
                           n17779, ZN => n10063);
   U3640 : OAI221_X1 port map( B1 => n1839, B2 => n19052, C1 => n5424, C2 => 
                           n19046, A => n9995, ZN => n9993);
   U3641 : AOI22_X1 port map( A1 => n19040, A2 => n17900, B1 => n19034, B2 => 
                           n17780, ZN => n9995);
   U3642 : OAI221_X1 port map( B1 => n1838, B2 => n19052, C1 => n5359, C2 => 
                           n19046, A => n9928, ZN => n9926);
   U3643 : AOI22_X1 port map( A1 => n19040, A2 => n17901, B1 => n19034, B2 => 
                           n17781, ZN => n9928);
   U3644 : OAI221_X1 port map( B1 => n1837, B2 => n19052, C1 => n5357, C2 => 
                           n19046, A => n9861, ZN => n9859);
   U3645 : AOI22_X1 port map( A1 => n19040, A2 => n17902, B1 => n19034, B2 => 
                           n17782, ZN => n9861);
   U3646 : OAI221_X1 port map( B1 => n1836, B2 => n19052, C1 => n5356, C2 => 
                           n19046, A => n9793, ZN => n9791);
   U3647 : AOI22_X1 port map( A1 => n19040, A2 => n17903, B1 => n19034, B2 => 
                           n17783, ZN => n9793);
   U3648 : OAI221_X1 port map( B1 => n1835, B2 => n19052, C1 => n5355, C2 => 
                           n19046, A => n9726, ZN => n9724);
   U3649 : AOI22_X1 port map( A1 => n19040, A2 => n17904, B1 => n19034, B2 => 
                           n17784, ZN => n9726);
   U3650 : OAI221_X1 port map( B1 => n1834, B2 => n19052, C1 => n5291, C2 => 
                           n19046, A => n9659, ZN => n9657);
   U3651 : AOI22_X1 port map( A1 => n19040, A2 => n17905, B1 => n19034, B2 => 
                           n17785, ZN => n9659);
   U3652 : OAI221_X1 port map( B1 => n1833, B2 => n19052, C1 => n5290, C2 => 
                           n19046, A => n9592, ZN => n9590);
   U3653 : AOI22_X1 port map( A1 => n19040, A2 => n17906, B1 => n19034, B2 => 
                           n17786, ZN => n9592);
   U3654 : OAI221_X1 port map( B1 => n1832, B2 => n19052, C1 => n5289, C2 => 
                           n19046, A => n9524, ZN => n9522);
   U3655 : AOI22_X1 port map( A1 => n19040, A2 => n17907, B1 => n19034, B2 => 
                           n17787, ZN => n9524);
   U3656 : OAI221_X1 port map( B1 => n1831, B2 => n19052, C1 => n5288, C2 => 
                           n19046, A => n9457, ZN => n9455);
   U3657 : AOI22_X1 port map( A1 => n19040, A2 => n17908, B1 => n19034, B2 => 
                           n17788, ZN => n9457);
   U3658 : OAI221_X1 port map( B1 => n1830, B2 => n19052, C1 => n5287, C2 => 
                           n19046, A => n9390, ZN => n9388);
   U3659 : AOI22_X1 port map( A1 => n19040, A2 => n17909, B1 => n19034, B2 => 
                           n17789, ZN => n9390);
   U3660 : OAI221_X1 port map( B1 => n1829, B2 => n19052, C1 => n5286, C2 => 
                           n19046, A => n9323, ZN => n9321);
   U3661 : AOI22_X1 port map( A1 => n19040, A2 => n17910, B1 => n19034, B2 => 
                           n17790, ZN => n9323);
   U3662 : OAI221_X1 port map( B1 => n1828, B2 => n19052, C1 => n5285, C2 => 
                           n19046, A => n7015, ZN => n7013);
   U3663 : AOI22_X1 port map( A1 => n19040, A2 => n17911, B1 => n19034, B2 => 
                           n17791, ZN => n7015);
   U3664 : OAI221_X1 port map( B1 => n4909, B2 => n19443, C1 => n2429, C2 => 
                           n19437, A => n10760, ZN => n10755);
   U3665 : AOI22_X1 port map( A1 => n19431, A2 => registers_4_12_port, B1 => 
                           n19425, B2 => n18004, ZN => n10760);
   U3666 : OAI221_X1 port map( B1 => n4908, B2 => n19443, C1 => n2428, C2 => 
                           n19437, A => n10692, ZN => n10687);
   U3667 : AOI22_X1 port map( A1 => n19431, A2 => registers_4_13_port, B1 => 
                           n19425, B2 => n18005, ZN => n10692);
   U3668 : OAI221_X1 port map( B1 => n4907, B2 => n19443, C1 => n2427, C2 => 
                           n19437, A => n10625, ZN => n10620);
   U3669 : AOI22_X1 port map( A1 => n19431, A2 => registers_4_14_port, B1 => 
                           n19425, B2 => n18006, ZN => n10625);
   U3670 : OAI221_X1 port map( B1 => n4906, B2 => n19443, C1 => n2426, C2 => 
                           n19437, A => n10558, ZN => n10553);
   U3671 : AOI22_X1 port map( A1 => n19431, A2 => registers_4_15_port, B1 => 
                           n19425, B2 => n18007, ZN => n10558);
   U3672 : OAI221_X1 port map( B1 => n4905, B2 => n19443, C1 => n2425, C2 => 
                           n19437, A => n10491, ZN => n10486);
   U3673 : AOI22_X1 port map( A1 => n19431, A2 => registers_4_16_port, B1 => 
                           n19425, B2 => n18008, ZN => n10491);
   U3674 : OAI221_X1 port map( B1 => n4904, B2 => n19443, C1 => n2424, C2 => 
                           n19437, A => n10423, ZN => n10418);
   U3675 : AOI22_X1 port map( A1 => n19431, A2 => registers_4_17_port, B1 => 
                           n19425, B2 => n18009, ZN => n10423);
   U3676 : OAI221_X1 port map( B1 => n4903, B2 => n19443, C1 => n2423, C2 => 
                           n19437, A => n10356, ZN => n10351);
   U3677 : AOI22_X1 port map( A1 => n19431, A2 => registers_4_18_port, B1 => 
                           n19425, B2 => n18010, ZN => n10356);
   U3678 : OAI221_X1 port map( B1 => n4902, B2 => n19443, C1 => n2422, C2 => 
                           n19437, A => n10289, ZN => n10284);
   U3679 : AOI22_X1 port map( A1 => n19431, A2 => registers_4_19_port, B1 => 
                           n19425, B2 => n18011, ZN => n10289);
   U3680 : OAI221_X1 port map( B1 => n4901, B2 => n19443, C1 => n2421, C2 => 
                           n19437, A => n10222, ZN => n10216);
   U3681 : AOI22_X1 port map( A1 => n19431, A2 => registers_4_20_port, B1 => 
                           n19425, B2 => n18012, ZN => n10222);
   U3682 : OAI221_X1 port map( B1 => n4900, B2 => n19443, C1 => n2420, C2 => 
                           n19437, A => n10154, ZN => n10149);
   U3683 : AOI22_X1 port map( A1 => n19431, A2 => registers_4_21_port, B1 => 
                           n19425, B2 => n18013, ZN => n10154);
   U3684 : OAI221_X1 port map( B1 => n4899, B2 => n19443, C1 => n2419, C2 => 
                           n19437, A => n10087, ZN => n10082);
   U3685 : AOI22_X1 port map( A1 => n19431, A2 => registers_4_22_port, B1 => 
                           n19425, B2 => n18014, ZN => n10087);
   U3686 : OAI221_X1 port map( B1 => n4898, B2 => n19443, C1 => n2418, C2 => 
                           n19437, A => n10020, ZN => n10015);
   U3687 : AOI22_X1 port map( A1 => n19431, A2 => registers_4_23_port, B1 => 
                           n19425, B2 => n18015, ZN => n10020);
   U3688 : OAI221_X1 port map( B1 => n4897, B2 => n19444, C1 => n2417, C2 => 
                           n19438, A => n9952, ZN => n9947);
   U3689 : AOI22_X1 port map( A1 => n19432, A2 => registers_4_24_port, B1 => 
                           n19426, B2 => n18016, ZN => n9952);
   U3690 : OAI221_X1 port map( B1 => n4896, B2 => n19444, C1 => n2416, C2 => 
                           n19438, A => n9885, ZN => n9880);
   U3691 : AOI22_X1 port map( A1 => n19432, A2 => registers_4_25_port, B1 => 
                           n19426, B2 => n18017, ZN => n9885);
   U3692 : OAI221_X1 port map( B1 => n4895, B2 => n19444, C1 => n2415, C2 => 
                           n19438, A => n9818, ZN => n9813);
   U3693 : AOI22_X1 port map( A1 => n19432, A2 => registers_4_26_port, B1 => 
                           n19426, B2 => n18018, ZN => n9818);
   U3694 : OAI221_X1 port map( B1 => n4894, B2 => n19444, C1 => n2414, C2 => 
                           n19438, A => n9751, ZN => n9746);
   U3695 : AOI22_X1 port map( A1 => n19432, A2 => registers_4_27_port, B1 => 
                           n19426, B2 => n18019, ZN => n9751);
   U3696 : OAI221_X1 port map( B1 => n4893, B2 => n19444, C1 => n2413, C2 => 
                           n19438, A => n9683, ZN => n9678);
   U3697 : AOI22_X1 port map( A1 => n19432, A2 => registers_4_28_port, B1 => 
                           n19426, B2 => n18020, ZN => n9683);
   U3698 : OAI221_X1 port map( B1 => n4892, B2 => n19444, C1 => n2412, C2 => 
                           n19438, A => n9616, ZN => n9611);
   U3699 : AOI22_X1 port map( A1 => n19432, A2 => registers_4_29_port, B1 => 
                           n19426, B2 => n18021, ZN => n9616);
   U3700 : OAI221_X1 port map( B1 => n4891, B2 => n19444, C1 => n2411, C2 => 
                           n19438, A => n9549, ZN => n9544);
   U3701 : AOI22_X1 port map( A1 => n19432, A2 => registers_4_30_port, B1 => 
                           n19426, B2 => n18022, ZN => n9549);
   U3702 : OAI221_X1 port map( B1 => n4890, B2 => n19444, C1 => n2410, C2 => 
                           n19438, A => n9482, ZN => n9476);
   U3703 : AOI22_X1 port map( A1 => n19432, A2 => registers_4_31_port, B1 => 
                           n19426, B2 => n18023, ZN => n9482);
   U3704 : OAI221_X1 port map( B1 => n4889, B2 => n19444, C1 => n2409, C2 => 
                           n19438, A => n9414, ZN => n9409);
   U3705 : AOI22_X1 port map( A1 => n19432, A2 => registers_4_32_port, B1 => 
                           n19426, B2 => n18024, ZN => n9414);
   U3706 : OAI221_X1 port map( B1 => n4888, B2 => n19444, C1 => n2408, C2 => 
                           n19438, A => n9347, ZN => n9342);
   U3707 : AOI22_X1 port map( A1 => n19432, A2 => registers_4_33_port, B1 => 
                           n19426, B2 => n18025, ZN => n9347);
   U3708 : OAI221_X1 port map( B1 => n4887, B2 => n19444, C1 => n2407, C2 => 
                           n19438, A => n9280, ZN => n9275);
   U3709 : AOI22_X1 port map( A1 => n19432, A2 => registers_4_34_port, B1 => 
                           n19426, B2 => n18026, ZN => n9280);
   U3710 : OAI221_X1 port map( B1 => n4886, B2 => n19444, C1 => n2406, C2 => 
                           n19438, A => n6973, ZN => n6968);
   U3711 : AOI22_X1 port map( A1 => n19432, A2 => registers_4_35_port, B1 => 
                           n19426, B2 => n18027, ZN => n6973);
   U3712 : OAI221_X1 port map( B1 => n4885, B2 => n19445, C1 => n2405, C2 => 
                           n19439, A => n6906, ZN => n6901);
   U3713 : AOI22_X1 port map( A1 => n19433, A2 => registers_4_36_port, B1 => 
                           n19427, B2 => n18028, ZN => n6906);
   U3714 : OAI221_X1 port map( B1 => n4884, B2 => n19445, C1 => n2404, C2 => 
                           n19439, A => n6839, ZN => n6834);
   U3715 : AOI22_X1 port map( A1 => n19433, A2 => registers_4_37_port, B1 => 
                           n19427, B2 => n18029, ZN => n6839);
   U3716 : OAI221_X1 port map( B1 => n4883, B2 => n19445, C1 => n2403, C2 => 
                           n19439, A => n6772, ZN => n6767);
   U3717 : AOI22_X1 port map( A1 => n19433, A2 => registers_4_38_port, B1 => 
                           n19427, B2 => n18030, ZN => n6772);
   U3718 : OAI221_X1 port map( B1 => n4882, B2 => n19445, C1 => n2402, C2 => 
                           n19439, A => n6705, ZN => n6700);
   U3719 : AOI22_X1 port map( A1 => n19433, A2 => registers_4_39_port, B1 => 
                           n19427, B2 => n18031, ZN => n6705);
   U3720 : OAI221_X1 port map( B1 => n4881, B2 => n19445, C1 => n2401, C2 => 
                           n19439, A => n6637, ZN => n6632);
   U3721 : AOI22_X1 port map( A1 => n19433, A2 => registers_4_40_port, B1 => 
                           n19427, B2 => n18032, ZN => n6637);
   U3722 : OAI221_X1 port map( B1 => n4880, B2 => n19445, C1 => n2400, C2 => 
                           n19439, A => n6571, ZN => n6566);
   U3723 : AOI22_X1 port map( A1 => n19433, A2 => registers_4_41_port, B1 => 
                           n19427, B2 => n18033, ZN => n6571);
   U3724 : OAI221_X1 port map( B1 => n4879, B2 => n19445, C1 => n2399, C2 => 
                           n19439, A => n6505, ZN => n6500);
   U3725 : AOI22_X1 port map( A1 => n19433, A2 => registers_4_42_port, B1 => 
                           n19427, B2 => n18034, ZN => n6505);
   U3726 : OAI221_X1 port map( B1 => n4878, B2 => n19445, C1 => n2398, C2 => 
                           n19439, A => n6439, ZN => n6434);
   U3727 : AOI22_X1 port map( A1 => n19433, A2 => registers_4_43_port, B1 => 
                           n19427, B2 => n18035, ZN => n6439);
   U3728 : OAI221_X1 port map( B1 => n4877, B2 => n19445, C1 => n2397, C2 => 
                           n19439, A => n6373, ZN => n6368);
   U3729 : AOI22_X1 port map( A1 => n19433, A2 => registers_4_44_port, B1 => 
                           n19427, B2 => n18036, ZN => n6373);
   U3730 : OAI221_X1 port map( B1 => n4876, B2 => n19445, C1 => n2396, C2 => 
                           n19439, A => n6307, ZN => n6302);
   U3731 : AOI22_X1 port map( A1 => n19433, A2 => registers_4_45_port, B1 => 
                           n19427, B2 => n18037, ZN => n6307);
   U3732 : OAI221_X1 port map( B1 => n4875, B2 => n19445, C1 => n2395, C2 => 
                           n19439, A => n6241, ZN => n6236);
   U3733 : AOI22_X1 port map( A1 => n19433, A2 => registers_4_46_port, B1 => 
                           n19427, B2 => n18038, ZN => n6241);
   U3734 : OAI221_X1 port map( B1 => n4874, B2 => n19445, C1 => n2394, C2 => 
                           n19439, A => n6175, ZN => n6170);
   U3735 : AOI22_X1 port map( A1 => n19433, A2 => registers_4_47_port, B1 => 
                           n19427, B2 => n18039, ZN => n6175);
   U3736 : OAI221_X1 port map( B1 => n4873, B2 => n19446, C1 => n2393, C2 => 
                           n19440, A => n6109, ZN => n6104);
   U3737 : AOI22_X1 port map( A1 => n19434, A2 => registers_4_48_port, B1 => 
                           n19428, B2 => n18040, ZN => n6109);
   U3738 : OAI221_X1 port map( B1 => n4872, B2 => n19446, C1 => n2392, C2 => 
                           n19440, A => n6043, ZN => n6038);
   U3739 : AOI22_X1 port map( A1 => n19434, A2 => registers_4_49_port, B1 => 
                           n19428, B2 => n18041, ZN => n6043);
   U3740 : OAI221_X1 port map( B1 => n4871, B2 => n19446, C1 => n2391, C2 => 
                           n19440, A => n5975, ZN => n5970);
   U3741 : AOI22_X1 port map( A1 => n19434, A2 => registers_4_50_port, B1 => 
                           n19428, B2 => n18042, ZN => n5975);
   U3742 : OAI221_X1 port map( B1 => n4870, B2 => n19446, C1 => n2390, C2 => 
                           n19440, A => n5907, ZN => n5902);
   U3743 : AOI22_X1 port map( A1 => n19434, A2 => registers_4_51_port, B1 => 
                           n19428, B2 => n18043, ZN => n5907);
   U3744 : OAI221_X1 port map( B1 => n4869, B2 => n19446, C1 => n2389, C2 => 
                           n19440, A => n5840, ZN => n5834);
   U3745 : AOI22_X1 port map( A1 => n19434, A2 => registers_4_52_port, B1 => 
                           n19428, B2 => n18044, ZN => n5840);
   U3746 : OAI221_X1 port map( B1 => n4868, B2 => n19446, C1 => n2388, C2 => 
                           n19440, A => n5773, ZN => n5762);
   U3747 : AOI22_X1 port map( A1 => n19434, A2 => registers_4_53_port, B1 => 
                           n19428, B2 => n18045, ZN => n5773);
   U3748 : OAI221_X1 port map( B1 => n4867, B2 => n19446, C1 => n2387, C2 => 
                           n19440, A => n5701, ZN => n5692);
   U3749 : AOI22_X1 port map( A1 => n19434, A2 => registers_4_54_port, B1 => 
                           n19428, B2 => n18046, ZN => n5701);
   U3750 : OAI221_X1 port map( B1 => n4866, B2 => n19446, C1 => n2386, C2 => 
                           n19440, A => n5631, ZN => n5624);
   U3751 : AOI22_X1 port map( A1 => n19434, A2 => registers_4_55_port, B1 => 
                           n19428, B2 => n18047, ZN => n5631);
   U3752 : OAI221_X1 port map( B1 => n4865, B2 => n19446, C1 => n2385, C2 => 
                           n19440, A => n5563, ZN => n5555);
   U3753 : AOI22_X1 port map( A1 => n19434, A2 => registers_4_56_port, B1 => 
                           n19428, B2 => n18048, ZN => n5563);
   U3754 : OAI221_X1 port map( B1 => n4864, B2 => n19446, C1 => n2384, C2 => 
                           n19440, A => n5493, ZN => n5486);
   U3755 : AOI22_X1 port map( A1 => n19434, A2 => registers_4_57_port, B1 => 
                           n19428, B2 => n18049, ZN => n5493);
   U3756 : OAI221_X1 port map( B1 => n4863, B2 => n19446, C1 => n2383, C2 => 
                           n19440, A => n5423, ZN => n5418);
   U3757 : AOI22_X1 port map( A1 => n19434, A2 => registers_4_58_port, B1 => 
                           n19428, B2 => n18050, ZN => n5423);
   U3758 : OAI221_X1 port map( B1 => n4862, B2 => n19446, C1 => n2382, C2 => 
                           n19440, A => n5353, ZN => n5348);
   U3759 : AOI22_X1 port map( A1 => n19434, A2 => registers_4_59_port, B1 => 
                           n19428, B2 => n18051, ZN => n5353);
   U3760 : OAI221_X1 port map( B1 => n1803, B2 => n19055, C1 => n5260, C2 => 
                           n19049, A => n5329, ZN => n5327);
   U3761 : AOI22_X1 port map( A1 => n19043, A2 => n17912, B1 => n19037, B2 => 
                           n17792, ZN => n5329);
   U3762 : OAI221_X1 port map( B1 => n1802, B2 => n19055, C1 => n5259, C2 => 
                           n19049, A => n4652, ZN => n4586);
   U3763 : AOI22_X1 port map( A1 => n19043, A2 => n17913, B1 => n19037, B2 => 
                           n17793, ZN => n4652);
   U3764 : OAI221_X1 port map( B1 => n1801, B2 => n19055, C1 => n5258, C2 => 
                           n19049, A => n3370, ZN => n3368);
   U3765 : AOI22_X1 port map( A1 => n19043, A2 => n17914, B1 => n19037, B2 => 
                           n17794, ZN => n3370);
   U3766 : OAI221_X1 port map( B1 => n1800, B2 => n19055, C1 => n5257, C2 => 
                           n19049, A => n3152, ZN => n3145);
   U3767 : AOI22_X1 port map( A1 => n19043, A2 => n17915, B1 => n19037, B2 => 
                           n17795, ZN => n3152);
   U3768 : OAI221_X1 port map( B1 => n1824, B2 => n19053, C1 => n5281, C2 => 
                           n19047, A => n6747, ZN => n6745);
   U3769 : AOI22_X1 port map( A1 => n19041, A2 => n17916, B1 => n19035, B2 => 
                           n17796, ZN => n6747);
   U3770 : OAI221_X1 port map( B1 => n1823, B2 => n19053, C1 => n5280, C2 => 
                           n19047, A => n6680, ZN => n6678);
   U3771 : AOI22_X1 port map( A1 => n19041, A2 => n17917, B1 => n19035, B2 => 
                           n17797, ZN => n6680);
   U3772 : OAI221_X1 port map( B1 => n1822, B2 => n19053, C1 => n5279, C2 => 
                           n19047, A => n6613, ZN => n6611);
   U3773 : AOI22_X1 port map( A1 => n19041, A2 => n17918, B1 => n19035, B2 => 
                           n17798, ZN => n6613);
   U3774 : OAI221_X1 port map( B1 => n1821, B2 => n19053, C1 => n5278, C2 => 
                           n19047, A => n6547, ZN => n6545);
   U3775 : AOI22_X1 port map( A1 => n19041, A2 => n17919, B1 => n19035, B2 => 
                           n17799, ZN => n6547);
   U3776 : OAI221_X1 port map( B1 => n1820, B2 => n19053, C1 => n5277, C2 => 
                           n19047, A => n6481, ZN => n6479);
   U3777 : AOI22_X1 port map( A1 => n19041, A2 => n17920, B1 => n19035, B2 => 
                           n17800, ZN => n6481);
   U3778 : OAI221_X1 port map( B1 => n1819, B2 => n19053, C1 => n5276, C2 => 
                           n19047, A => n6415, ZN => n6413);
   U3779 : AOI22_X1 port map( A1 => n19041, A2 => n17921, B1 => n19035, B2 => 
                           n17801, ZN => n6415);
   U3780 : OAI221_X1 port map( B1 => n1818, B2 => n19053, C1 => n5275, C2 => 
                           n19047, A => n6349, ZN => n6347);
   U3781 : AOI22_X1 port map( A1 => n19041, A2 => n17922, B1 => n19035, B2 => 
                           n17802, ZN => n6349);
   U3782 : OAI221_X1 port map( B1 => n1817, B2 => n19053, C1 => n5274, C2 => 
                           n19047, A => n6283, ZN => n6281);
   U3783 : AOI22_X1 port map( A1 => n19041, A2 => n17923, B1 => n19035, B2 => 
                           n17803, ZN => n6283);
   U3784 : OAI221_X1 port map( B1 => n1816, B2 => n19053, C1 => n5273, C2 => 
                           n19047, A => n6217, ZN => n6215);
   U3785 : AOI22_X1 port map( A1 => n19041, A2 => n17924, B1 => n19035, B2 => 
                           n17804, ZN => n6217);
   U3786 : OAI221_X1 port map( B1 => n1827, B2 => n19053, C1 => n5284, C2 => 
                           n19047, A => n6949, ZN => n6947);
   U3787 : AOI22_X1 port map( A1 => n19041, A2 => n17925, B1 => n19035, B2 => 
                           n17805, ZN => n6949);
   U3788 : OAI221_X1 port map( B1 => n1826, B2 => n19053, C1 => n5283, C2 => 
                           n19047, A => n6882, ZN => n6880);
   U3789 : AOI22_X1 port map( A1 => n19041, A2 => n17926, B1 => n19035, B2 => 
                           n17806, ZN => n6882);
   U3790 : OAI221_X1 port map( B1 => n4921, B2 => n19442, C1 => n2441, C2 => 
                           n19436, A => n11592, ZN => n11582);
   U3791 : AOI22_X1 port map( A1 => n19430, A2 => registers_4_0_port, B1 => 
                           n19424, B2 => n11593, ZN => n11592);
   U3792 : OAI221_X1 port map( B1 => n4920, B2 => n19442, C1 => n2440, C2 => 
                           n19436, A => n11500, ZN => n11495);
   U3793 : AOI22_X1 port map( A1 => n19430, A2 => registers_4_1_port, B1 => 
                           n19424, B2 => n11501, ZN => n11500);
   U3794 : OAI221_X1 port map( B1 => n4919, B2 => n19442, C1 => n2439, C2 => 
                           n19436, A => n11432, ZN => n11427);
   U3795 : AOI22_X1 port map( A1 => n19430, A2 => registers_4_2_port, B1 => 
                           n19424, B2 => n11433, ZN => n11432);
   U3796 : OAI221_X1 port map( B1 => n4918, B2 => n19442, C1 => n2438, C2 => 
                           n19436, A => n11365, ZN => n11360);
   U3797 : AOI22_X1 port map( A1 => n19430, A2 => registers_4_3_port, B1 => 
                           n19424, B2 => n11366, ZN => n11365);
   U3798 : OAI221_X1 port map( B1 => n4917, B2 => n19442, C1 => n2437, C2 => 
                           n19436, A => n11298, ZN => n11293);
   U3799 : AOI22_X1 port map( A1 => n19430, A2 => registers_4_4_port, B1 => 
                           n19424, B2 => n17996, ZN => n11298);
   U3800 : OAI221_X1 port map( B1 => n4916, B2 => n19442, C1 => n2436, C2 => 
                           n19436, A => n11231, ZN => n11226);
   U3801 : AOI22_X1 port map( A1 => n19430, A2 => registers_4_5_port, B1 => 
                           n19424, B2 => n17997, ZN => n11231);
   U3802 : OAI221_X1 port map( B1 => n4915, B2 => n19442, C1 => n2435, C2 => 
                           n19436, A => n11163, ZN => n11158);
   U3803 : AOI22_X1 port map( A1 => n19430, A2 => registers_4_6_port, B1 => 
                           n19424, B2 => n17998, ZN => n11163);
   U3804 : OAI221_X1 port map( B1 => n4914, B2 => n19442, C1 => n2434, C2 => 
                           n19436, A => n11096, ZN => n11091);
   U3805 : AOI22_X1 port map( A1 => n19430, A2 => registers_4_7_port, B1 => 
                           n19424, B2 => n17999, ZN => n11096);
   U3806 : OAI221_X1 port map( B1 => n4913, B2 => n19442, C1 => n2433, C2 => 
                           n19436, A => n11029, ZN => n11024);
   U3807 : AOI22_X1 port map( A1 => n19430, A2 => registers_4_8_port, B1 => 
                           n19424, B2 => n18000, ZN => n11029);
   U3808 : OAI221_X1 port map( B1 => n4912, B2 => n19442, C1 => n2432, C2 => 
                           n19436, A => n10962, ZN => n10956);
   U3809 : AOI22_X1 port map( A1 => n19430, A2 => registers_4_9_port, B1 => 
                           n19424, B2 => n18001, ZN => n10962);
   U3810 : OAI221_X1 port map( B1 => n4911, B2 => n19442, C1 => n2431, C2 => 
                           n19436, A => n10894, ZN => n10889);
   U3811 : AOI22_X1 port map( A1 => n19430, A2 => registers_4_10_port, B1 => 
                           n19424, B2 => n18002, ZN => n10894);
   U3812 : OAI221_X1 port map( B1 => n4910, B2 => n19442, C1 => n2430, C2 => 
                           n19436, A => n10827, ZN => n10822);
   U3813 : AOI22_X1 port map( A1 => n19430, A2 => registers_4_11_port, B1 => 
                           n19424, B2 => n18003, ZN => n10827);
   U3814 : OAI221_X1 port map( B1 => n1863, B2 => n19050, C1 => n6033, C2 => 
                           n19044, A => n11678, ZN => n11668);
   U3815 : AOI22_X1 port map( A1 => n19038, A2 => n11606, B1 => n19032, B2 => 
                           n11586, ZN => n11678);
   U3816 : OAI221_X1 port map( B1 => n1862, B2 => n19050, C1 => n5968, C2 => 
                           n19044, A => n11543, ZN => n11540);
   U3817 : AOI22_X1 port map( A1 => n19038, A2 => n11507, B1 => n19032, B2 => 
                           n11499, ZN => n11543);
   U3818 : OAI221_X1 port map( B1 => n1861, B2 => n19050, C1 => n5966, C2 => 
                           n19044, A => n11475, ZN => n11473);
   U3819 : AOI22_X1 port map( A1 => n19038, A2 => n11440, B1 => n19032, B2 => 
                           n11431, ZN => n11475);
   U3820 : OAI221_X1 port map( B1 => n1860, B2 => n19050, C1 => n5901, C2 => 
                           n19044, A => n11408, ZN => n11406);
   U3821 : AOI22_X1 port map( A1 => n19038, A2 => n11372, B1 => n19032, B2 => 
                           n11364, ZN => n11408);
   U3822 : OAI221_X1 port map( B1 => n1859, B2 => n19050, C1 => n5835, C2 => 
                           n19044, A => n11341, ZN => n11339);
   U3823 : AOI22_X1 port map( A1 => n19038, A2 => n17927, B1 => n19032, B2 => 
                           n17807, ZN => n11341);
   U3824 : OAI221_X1 port map( B1 => n1858, B2 => n19050, C1 => n5769, C2 => 
                           n19044, A => n11273, ZN => n11271);
   U3825 : AOI22_X1 port map( A1 => n19038, A2 => n17928, B1 => n19032, B2 => 
                           n17808, ZN => n11273);
   U3826 : OAI221_X1 port map( B1 => n1857, B2 => n19050, C1 => n5767, C2 => 
                           n19044, A => n11206, ZN => n11204);
   U3827 : AOI22_X1 port map( A1 => n19038, A2 => n17929, B1 => n19032, B2 => 
                           n17809, ZN => n11206);
   U3828 : OAI221_X1 port map( B1 => n1856, B2 => n19050, C1 => n5766, C2 => 
                           n19044, A => n11139, ZN => n11137);
   U3829 : AOI22_X1 port map( A1 => n19038, A2 => n17930, B1 => n19032, B2 => 
                           n17810, ZN => n11139);
   U3830 : OAI221_X1 port map( B1 => n1855, B2 => n19050, C1 => n5765, C2 => 
                           n19044, A => n11072, ZN => n11070);
   U3831 : AOI22_X1 port map( A1 => n19038, A2 => n17931, B1 => n19032, B2 => 
                           n17811, ZN => n11072);
   U3832 : OAI221_X1 port map( B1 => n1854, B2 => n19050, C1 => n5764, C2 => 
                           n19044, A => n11004, ZN => n11002);
   U3833 : AOI22_X1 port map( A1 => n19038, A2 => n17932, B1 => n19032, B2 => 
                           n17812, ZN => n11004);
   U3834 : OAI221_X1 port map( B1 => n1853, B2 => n19050, C1 => n5763, C2 => 
                           n19044, A => n10937, ZN => n10935);
   U3835 : AOI22_X1 port map( A1 => n19038, A2 => n17933, B1 => n19032, B2 => 
                           n17813, ZN => n10937);
   U3836 : OAI221_X1 port map( B1 => n1852, B2 => n19050, C1 => n5698, C2 => 
                           n19044, A => n10870, ZN => n10868);
   U3837 : AOI22_X1 port map( A1 => n19038, A2 => n17934, B1 => n19032, B2 => 
                           n17814, ZN => n10870);
   U3838 : OAI221_X1 port map( B1 => n3354, B2 => n19220, C1 => n4838, C2 => 
                           n19214, A => n10786, ZN => n10781);
   U3839 : AOI22_X1 port map( A1 => n19208, A2 => n17816, B1 => n19202, B2 => 
                           n18056, ZN => n10786);
   U3840 : OAI221_X1 port map( B1 => n3353, B2 => n19220, C1 => n4837, C2 => 
                           n19214, A => n10719, ZN => n10714);
   U3841 : AOI22_X1 port map( A1 => n19208, A2 => n17817, B1 => n19202, B2 => 
                           n18057, ZN => n10719);
   U3842 : OAI221_X1 port map( B1 => n3352, B2 => n19220, C1 => n4836, C2 => 
                           n19214, A => n10652, ZN => n10647);
   U3843 : AOI22_X1 port map( A1 => n19208, A2 => n17818, B1 => n19202, B2 => 
                           n18058, ZN => n10652);
   U3844 : OAI221_X1 port map( B1 => n3351, B2 => n19220, C1 => n4835, C2 => 
                           n19214, A => n10584, ZN => n10579);
   U3845 : AOI22_X1 port map( A1 => n19208, A2 => n17819, B1 => n19202, B2 => 
                           n18059, ZN => n10584);
   U3846 : OAI221_X1 port map( B1 => n3350, B2 => n19220, C1 => n4834, C2 => 
                           n19214, A => n10517, ZN => n10512);
   U3847 : AOI22_X1 port map( A1 => n19208, A2 => n17820, B1 => n19202, B2 => 
                           n18060, ZN => n10517);
   U3848 : OAI221_X1 port map( B1 => n3349, B2 => n19220, C1 => n4833, C2 => 
                           n19214, A => n10450, ZN => n10445);
   U3849 : AOI22_X1 port map( A1 => n19208, A2 => n17821, B1 => n19202, B2 => 
                           n18061, ZN => n10450);
   U3850 : OAI221_X1 port map( B1 => n3348, B2 => n19220, C1 => n4832, C2 => 
                           n19214, A => n10383, ZN => n10378);
   U3851 : AOI22_X1 port map( A1 => n19208, A2 => n17822, B1 => n19202, B2 => 
                           n18062, ZN => n10383);
   U3852 : OAI221_X1 port map( B1 => n3347, B2 => n19220, C1 => n4831, C2 => 
                           n19214, A => n10315, ZN => n10310);
   U3853 : AOI22_X1 port map( A1 => n19208, A2 => n17823, B1 => n19202, B2 => 
                           n18063, ZN => n10315);
   U3854 : OAI221_X1 port map( B1 => n3346, B2 => n19220, C1 => n4830, C2 => 
                           n19214, A => n10248, ZN => n10243);
   U3855 : AOI22_X1 port map( A1 => n19208, A2 => n17824, B1 => n19202, B2 => 
                           n18064, ZN => n10248);
   U3856 : OAI221_X1 port map( B1 => n3345, B2 => n19220, C1 => n4829, C2 => 
                           n19214, A => n10181, ZN => n10176);
   U3857 : AOI22_X1 port map( A1 => n19208, A2 => n17825, B1 => n19202, B2 => 
                           n18065, ZN => n10181);
   U3858 : OAI221_X1 port map( B1 => n3344, B2 => n19220, C1 => n4828, C2 => 
                           n19214, A => n10114, ZN => n10108);
   U3859 : AOI22_X1 port map( A1 => n19208, A2 => n17826, B1 => n19202, B2 => 
                           n18066, ZN => n10114);
   U3860 : OAI221_X1 port map( B1 => n3343, B2 => n19220, C1 => n4827, C2 => 
                           n19214, A => n10046, ZN => n10041);
   U3861 : AOI22_X1 port map( A1 => n19208, A2 => n17827, B1 => n19202, B2 => 
                           n18067, ZN => n10046);
   U3862 : OAI221_X1 port map( B1 => n3342, B2 => n19221, C1 => n4826, C2 => 
                           n19215, A => n9979, ZN => n9974);
   U3863 : AOI22_X1 port map( A1 => n19209, A2 => n17828, B1 => n19203, B2 => 
                           n18068, ZN => n9979);
   U3864 : OAI221_X1 port map( B1 => n3341, B2 => n19221, C1 => n4825, C2 => 
                           n19215, A => n9912, ZN => n9907);
   U3865 : AOI22_X1 port map( A1 => n19209, A2 => n17829, B1 => n19203, B2 => 
                           n18069, ZN => n9912);
   U3866 : OAI221_X1 port map( B1 => n3340, B2 => n19221, C1 => n4824, C2 => 
                           n19215, A => n9844, ZN => n9839);
   U3867 : AOI22_X1 port map( A1 => n19209, A2 => n17830, B1 => n19203, B2 => 
                           n18070, ZN => n9844);
   U3868 : OAI221_X1 port map( B1 => n3339, B2 => n19221, C1 => n4823, C2 => 
                           n19215, A => n9777, ZN => n9772);
   U3869 : AOI22_X1 port map( A1 => n19209, A2 => n17831, B1 => n19203, B2 => 
                           n18071, ZN => n9777);
   U3870 : OAI221_X1 port map( B1 => n3338, B2 => n19221, C1 => n4822, C2 => 
                           n19215, A => n9710, ZN => n9705);
   U3871 : AOI22_X1 port map( A1 => n19209, A2 => n17832, B1 => n19203, B2 => 
                           n18072, ZN => n9710);
   U3872 : OAI221_X1 port map( B1 => n3337, B2 => n19221, C1 => n4821, C2 => 
                           n19215, A => n9643, ZN => n9638);
   U3873 : AOI22_X1 port map( A1 => n19209, A2 => n17833, B1 => n19203, B2 => 
                           n18073, ZN => n9643);
   U3874 : OAI221_X1 port map( B1 => n3336, B2 => n19221, C1 => n4820, C2 => 
                           n19215, A => n9575, ZN => n9570);
   U3875 : AOI22_X1 port map( A1 => n19209, A2 => n17834, B1 => n19203, B2 => 
                           n18074, ZN => n9575);
   U3876 : OAI221_X1 port map( B1 => n3335, B2 => n19221, C1 => n4819, C2 => 
                           n19215, A => n9508, ZN => n9503);
   U3877 : AOI22_X1 port map( A1 => n19209, A2 => n17835, B1 => n19203, B2 => 
                           n18075, ZN => n9508);
   U3878 : OAI221_X1 port map( B1 => n3334, B2 => n19221, C1 => n4818, C2 => 
                           n19215, A => n9441, ZN => n9436);
   U3879 : AOI22_X1 port map( A1 => n19209, A2 => n17836, B1 => n19203, B2 => 
                           n18076, ZN => n9441);
   U3880 : OAI221_X1 port map( B1 => n3333, B2 => n19221, C1 => n4817, C2 => 
                           n19215, A => n9374, ZN => n9368);
   U3881 : AOI22_X1 port map( A1 => n19209, A2 => n17837, B1 => n19203, B2 => 
                           n18077, ZN => n9374);
   U3882 : OAI221_X1 port map( B1 => n3332, B2 => n19221, C1 => n4816, C2 => 
                           n19215, A => n9306, ZN => n9301);
   U3883 : AOI22_X1 port map( A1 => n19209, A2 => n17838, B1 => n19203, B2 => 
                           n18078, ZN => n9306);
   U3884 : OAI221_X1 port map( B1 => n3331, B2 => n19221, C1 => n4815, C2 => 
                           n19215, A => n6999, ZN => n6994);
   U3885 : AOI22_X1 port map( A1 => n19209, A2 => n17839, B1 => n19203, B2 => 
                           n18079, ZN => n6999);
   U3886 : OAI221_X1 port map( B1 => n3330, B2 => n19222, C1 => n4814, C2 => 
                           n19216, A => n6932, ZN => n6927);
   U3887 : AOI22_X1 port map( A1 => n19210, A2 => n17840, B1 => n19204, B2 => 
                           n18080, ZN => n6932);
   U3888 : OAI221_X1 port map( B1 => n3329, B2 => n19222, C1 => n4813, C2 => 
                           n19216, A => n6865, ZN => n6860);
   U3889 : AOI22_X1 port map( A1 => n19210, A2 => n17841, B1 => n19204, B2 => 
                           n18081, ZN => n6865);
   U3890 : OAI221_X1 port map( B1 => n3328, B2 => n19222, C1 => n4812, C2 => 
                           n19216, A => n6798, ZN => n6793);
   U3891 : AOI22_X1 port map( A1 => n19210, A2 => n17842, B1 => n19204, B2 => 
                           n18082, ZN => n6798);
   U3892 : OAI221_X1 port map( B1 => n3327, B2 => n19222, C1 => n4811, C2 => 
                           n19216, A => n6731, ZN => n6726);
   U3893 : AOI22_X1 port map( A1 => n19210, A2 => n17843, B1 => n19204, B2 => 
                           n18083, ZN => n6731);
   U3894 : OAI221_X1 port map( B1 => n3326, B2 => n19222, C1 => n4810, C2 => 
                           n19216, A => n6664, ZN => n6659);
   U3895 : AOI22_X1 port map( A1 => n19210, A2 => n17844, B1 => n19204, B2 => 
                           n18084, ZN => n6664);
   U3896 : OAI221_X1 port map( B1 => n3325, B2 => n19222, C1 => n4809, C2 => 
                           n19216, A => n6597, ZN => n6592);
   U3897 : AOI22_X1 port map( A1 => n19210, A2 => n17845, B1 => n19204, B2 => 
                           n18085, ZN => n6597);
   U3898 : OAI221_X1 port map( B1 => n3324, B2 => n19222, C1 => n4808, C2 => 
                           n19216, A => n6531, ZN => n6526);
   U3899 : AOI22_X1 port map( A1 => n19210, A2 => n17846, B1 => n19204, B2 => 
                           n18086, ZN => n6531);
   U3900 : OAI221_X1 port map( B1 => n3323, B2 => n19222, C1 => n4807, C2 => 
                           n19216, A => n6465, ZN => n6460);
   U3901 : AOI22_X1 port map( A1 => n19210, A2 => n17847, B1 => n19204, B2 => 
                           n18087, ZN => n6465);
   U3902 : OAI221_X1 port map( B1 => n3322, B2 => n19222, C1 => n4806, C2 => 
                           n19216, A => n6399, ZN => n6394);
   U3903 : AOI22_X1 port map( A1 => n19210, A2 => n17848, B1 => n19204, B2 => 
                           n18088, ZN => n6399);
   U3904 : OAI221_X1 port map( B1 => n3321, B2 => n19222, C1 => n4805, C2 => 
                           n19216, A => n6333, ZN => n6328);
   U3905 : AOI22_X1 port map( A1 => n19210, A2 => n17849, B1 => n19204, B2 => 
                           n18089, ZN => n6333);
   U3906 : OAI221_X1 port map( B1 => n3320, B2 => n19222, C1 => n4804, C2 => 
                           n19216, A => n6267, ZN => n6262);
   U3907 : AOI22_X1 port map( A1 => n19210, A2 => n17850, B1 => n19204, B2 => 
                           n18090, ZN => n6267);
   U3908 : OAI221_X1 port map( B1 => n3319, B2 => n19222, C1 => n4803, C2 => 
                           n19216, A => n6201, ZN => n6196);
   U3909 : AOI22_X1 port map( A1 => n19210, A2 => n17851, B1 => n19204, B2 => 
                           n18091, ZN => n6201);
   U3910 : OAI221_X1 port map( B1 => n3318, B2 => n19223, C1 => n4802, C2 => 
                           n19217, A => n6135, ZN => n6130);
   U3911 : AOI22_X1 port map( A1 => n19211, A2 => n17852, B1 => n19205, B2 => 
                           n18092, ZN => n6135);
   U3912 : OAI221_X1 port map( B1 => n3317, B2 => n19223, C1 => n4801, C2 => 
                           n19217, A => n6069, ZN => n6064);
   U3913 : AOI22_X1 port map( A1 => n19211, A2 => n17853, B1 => n19205, B2 => 
                           n18093, ZN => n6069);
   U3914 : OAI221_X1 port map( B1 => n3316, B2 => n19223, C1 => n4800, C2 => 
                           n19217, A => n6001, ZN => n5996);
   U3915 : AOI22_X1 port map( A1 => n19211, A2 => n17854, B1 => n19205, B2 => 
                           n18094, ZN => n6001);
   U3916 : OAI221_X1 port map( B1 => n3315, B2 => n19223, C1 => n4799, C2 => 
                           n19217, A => n5933, ZN => n5928);
   U3917 : AOI22_X1 port map( A1 => n19211, A2 => n17855, B1 => n19205, B2 => 
                           n18095, ZN => n5933);
   U3918 : OAI221_X1 port map( B1 => n3314, B2 => n19223, C1 => n4798, C2 => 
                           n19217, A => n5866, ZN => n5861);
   U3919 : AOI22_X1 port map( A1 => n19211, A2 => n17856, B1 => n19205, B2 => 
                           n18096, ZN => n5866);
   U3920 : OAI221_X1 port map( B1 => n3313, B2 => n19223, C1 => n4797, C2 => 
                           n19217, A => n5799, ZN => n5794);
   U3921 : AOI22_X1 port map( A1 => n19211, A2 => n17857, B1 => n19205, B2 => 
                           n18097, ZN => n5799);
   U3922 : OAI221_X1 port map( B1 => n3312, B2 => n19223, C1 => n4796, C2 => 
                           n19217, A => n5727, ZN => n5722);
   U3923 : AOI22_X1 port map( A1 => n19211, A2 => n17858, B1 => n19205, B2 => 
                           n18098, ZN => n5727);
   U3924 : OAI221_X1 port map( B1 => n3311, B2 => n19223, C1 => n4795, C2 => 
                           n19217, A => n5657, ZN => n5652);
   U3925 : AOI22_X1 port map( A1 => n19211, A2 => n17859, B1 => n19205, B2 => 
                           n18099, ZN => n5657);
   U3926 : OAI221_X1 port map( B1 => n3310, B2 => n19223, C1 => n4794, C2 => 
                           n19217, A => n5589, ZN => n5584);
   U3927 : AOI22_X1 port map( A1 => n19211, A2 => n17860, B1 => n19205, B2 => 
                           n18100, ZN => n5589);
   U3928 : OAI221_X1 port map( B1 => n3309, B2 => n19223, C1 => n4793, C2 => 
                           n19217, A => n5520, ZN => n5515);
   U3929 : AOI22_X1 port map( A1 => n19211, A2 => n17861, B1 => n19205, B2 => 
                           n18101, ZN => n5520);
   U3930 : OAI221_X1 port map( B1 => n3308, B2 => n19223, C1 => n4792, C2 => 
                           n19217, A => n5451, ZN => n5446);
   U3931 : AOI22_X1 port map( A1 => n19211, A2 => n17862, B1 => n19205, B2 => 
                           n18102, ZN => n5451);
   U3932 : OAI221_X1 port map( B1 => n3307, B2 => n19223, C1 => n4791, C2 => 
                           n19217, A => n5383, ZN => n5378);
   U3933 : AOI22_X1 port map( A1 => n19211, A2 => n17863, B1 => n19205, B2 => 
                           n18103, ZN => n5383);
   U3934 : OAI221_X1 port map( B1 => n3306, B2 => n19224, C1 => n4790, C2 => 
                           n19218, A => n5313, ZN => n5308);
   U3935 : AOI22_X1 port map( A1 => n19212, A2 => n17864, B1 => n19206, B2 => 
                           n18104, ZN => n5313);
   U3936 : OAI221_X1 port map( B1 => n3306, B2 => n19423, C1 => n4790, C2 => 
                           n19417, A => n5254, ZN => n5054);
   U3937 : AOI22_X1 port map( A1 => n19411, A2 => n17864, B1 => n19405, B2 => 
                           n18104, ZN => n5254);
   U3938 : OAI221_X1 port map( B1 => n3305, B2 => n19224, C1 => n4789, C2 => 
                           n19218, A => n4380, ZN => n4311);
   U3939 : AOI22_X1 port map( A1 => n19212, A2 => n17865, B1 => n19206, B2 => 
                           n18105, ZN => n4380);
   U3940 : OAI221_X1 port map( B1 => n3305, B2 => n19423, C1 => n4789, C2 => 
                           n19417, A => n3972, ZN => n3772);
   U3941 : AOI22_X1 port map( A1 => n19411, A2 => n17865, B1 => n19405, B2 => 
                           n18105, ZN => n3972);
   U3942 : OAI221_X1 port map( B1 => n3304, B2 => n19224, C1 => n4788, C2 => 
                           n19218, A => n3284, ZN => n3274);
   U3943 : AOI22_X1 port map( A1 => n19212, A2 => n17866, B1 => n19206, B2 => 
                           n18106, ZN => n3284);
   U3944 : OAI221_X1 port map( B1 => n3304, B2 => n19423, C1 => n4788, C2 => 
                           n19417, A => n3236, ZN => n3220);
   U3945 : AOI22_X1 port map( A1 => n19411, A2 => n17866, B1 => n19405, B2 => 
                           n18106, ZN => n3236);
   U3946 : OAI221_X1 port map( B1 => n3303, B2 => n19224, C1 => n4787, C2 => 
                           n19218, A => n3108, ZN => n3029);
   U3947 : AOI22_X1 port map( A1 => n19212, A2 => n17867, B1 => n19206, B2 => 
                           n18107, ZN => n3108);
   U3948 : OAI221_X1 port map( B1 => n3303, B2 => n19423, C1 => n4787, C2 => 
                           n19417, A => n2987, ZN => n2777);
   U3949 : AOI22_X1 port map( A1 => n19411, A2 => n17867, B1 => n19405, B2 => 
                           n18107, ZN => n2987);
   U3950 : OAI221_X1 port map( B1 => n3366, B2 => n19219, C1 => n4850, C2 => 
                           n19213, A => n11641, ZN => n11629);
   U3951 : AOI22_X1 port map( A1 => n19207, A2 => n11598, B1 => n19201, B2 => 
                           n11599, ZN => n11641);
   U3952 : OAI221_X1 port map( B1 => n3365, B2 => n19219, C1 => n4849, C2 => 
                           n19213, A => n11526, ZN => n11521);
   U3953 : AOI22_X1 port map( A1 => n19207, A2 => n11503, B1 => n19201, B2 => 
                           n11504, ZN => n11526);
   U3954 : OAI221_X1 port map( B1 => n3364, B2 => n19219, C1 => n4848, C2 => 
                           n19213, A => n11459, ZN => n11454);
   U3955 : AOI22_X1 port map( A1 => n19207, A2 => n11435, B1 => n19201, B2 => 
                           n11437, ZN => n11459);
   U3956 : OAI221_X1 port map( B1 => n3363, B2 => n19219, C1 => n4847, C2 => 
                           n19213, A => n11392, ZN => n11387);
   U3957 : AOI22_X1 port map( A1 => n19207, A2 => n11368, B1 => n19201, B2 => 
                           n11369, ZN => n11392);
   U3958 : OAI221_X1 port map( B1 => n3362, B2 => n19219, C1 => n4846, C2 => 
                           n19213, A => n11324, ZN => n11319);
   U3959 : AOI22_X1 port map( A1 => n19207, A2 => n17868, B1 => n19201, B2 => 
                           n18108, ZN => n11324);
   U3960 : OAI221_X1 port map( B1 => n3361, B2 => n19219, C1 => n4845, C2 => 
                           n19213, A => n11257, ZN => n11252);
   U3961 : AOI22_X1 port map( A1 => n19207, A2 => n17869, B1 => n19201, B2 => 
                           n18109, ZN => n11257);
   U3962 : OAI221_X1 port map( B1 => n3360, B2 => n19219, C1 => n4844, C2 => 
                           n19213, A => n11190, ZN => n11185);
   U3963 : AOI22_X1 port map( A1 => n19207, A2 => n17870, B1 => n19201, B2 => 
                           n18110, ZN => n11190);
   U3964 : OAI221_X1 port map( B1 => n3359, B2 => n19219, C1 => n4843, C2 => 
                           n19213, A => n11123, ZN => n11117);
   U3965 : AOI22_X1 port map( A1 => n19207, A2 => n17871, B1 => n19201, B2 => 
                           n18111, ZN => n11123);
   U3966 : OAI221_X1 port map( B1 => n3358, B2 => n19219, C1 => n4842, C2 => 
                           n19213, A => n11055, ZN => n11050);
   U3967 : AOI22_X1 port map( A1 => n19207, A2 => n17872, B1 => n19201, B2 => 
                           n18112, ZN => n11055);
   U3968 : OAI221_X1 port map( B1 => n3357, B2 => n19219, C1 => n4841, C2 => 
                           n19213, A => n10988, ZN => n10983);
   U3969 : AOI22_X1 port map( A1 => n19207, A2 => n17873, B1 => n19201, B2 => 
                           n18113, ZN => n10988);
   U3970 : OAI221_X1 port map( B1 => n3356, B2 => n19219, C1 => n4840, C2 => 
                           n19213, A => n10921, ZN => n10916);
   U3971 : AOI22_X1 port map( A1 => n19207, A2 => n17874, B1 => n19201, B2 => 
                           n18114, ZN => n10921);
   U3972 : OAI221_X1 port map( B1 => n3355, B2 => n19219, C1 => n4839, C2 => 
                           n19213, A => n10853, ZN => n10848);
   U3973 : AOI22_X1 port map( A1 => n19207, A2 => n17875, B1 => n19201, B2 => 
                           n18115, ZN => n10853);
   U3974 : AOI22_X1 port map( A1 => n19041, A2 => n17935, B1 => n19035, B2 => 
                           n17815, ZN => n6815);
   U3975 : OAI221_X1 port map( B1 => n3577, B2 => n18965, C1 => n18959, C2 => 
                           n2447, A => n5335, ZN => n5333);
   U3976 : AOI22_X1 port map( A1 => n18953, A2 => n18117, B1 => n18947, B2 => 
                           n17697, ZN => n5335);
   U3977 : OAI221_X1 port map( B1 => n3576, B2 => n18965, C1 => n18959, C2 => 
                           n2446, A => n4786, ZN => n4784);
   U3978 : AOI22_X1 port map( A1 => n18953, A2 => n18118, B1 => n18947, B2 => 
                           n17698, ZN => n4786);
   U3979 : OAI221_X1 port map( B1 => n3575, B2 => n18965, C1 => n18959, C2 => 
                           n2445, A => n3504, ZN => n3438);
   U3980 : AOI22_X1 port map( A1 => n18953, A2 => n18119, B1 => n18947, B2 => 
                           n17699, ZN => n3504);
   U3981 : OAI221_X1 port map( B1 => n3574, B2 => n18965, C1 => n18959, C2 => 
                           n2444, A => n3178, ZN => n3167);
   U3982 : AOI22_X1 port map( A1 => n18953, A2 => n18120, B1 => n18947, B2 => 
                           n17700, ZN => n3178);
   U3983 : OAI221_X1 port map( B1 => n3598, B2 => n18963, C1 => n18957, C2 => 
                           n2724, A => n6754, ZN => n6752);
   U3984 : AOI22_X1 port map( A1 => n18951, A2 => n18121, B1 => n18945, B2 => 
                           n17701, ZN => n6754);
   U3985 : OAI221_X1 port map( B1 => n3597, B2 => n18963, C1 => n18957, C2 => 
                           n2723, A => n6686, ZN => n6684);
   U3986 : AOI22_X1 port map( A1 => n18951, A2 => n18122, B1 => n18945, B2 => 
                           n17702, ZN => n6686);
   U3987 : OAI221_X1 port map( B1 => n3596, B2 => n18963, C1 => n18957, C2 => 
                           n2722, A => n6619, ZN => n6617);
   U3988 : AOI22_X1 port map( A1 => n18951, A2 => n18123, B1 => n18945, B2 => 
                           n17703, ZN => n6619);
   U3989 : OAI221_X1 port map( B1 => n3595, B2 => n18963, C1 => n18957, C2 => 
                           n2721, A => n6553, ZN => n6551);
   U3990 : AOI22_X1 port map( A1 => n18951, A2 => n18124, B1 => n18945, B2 => 
                           n17704, ZN => n6553);
   U3991 : OAI221_X1 port map( B1 => n3594, B2 => n18963, C1 => n18957, C2 => 
                           n2720, A => n6487, ZN => n6485);
   U3992 : AOI22_X1 port map( A1 => n18951, A2 => n18125, B1 => n18945, B2 => 
                           n17705, ZN => n6487);
   U3993 : OAI221_X1 port map( B1 => n3593, B2 => n18963, C1 => n18957, C2 => 
                           n2463, A => n6421, ZN => n6419);
   U3994 : AOI22_X1 port map( A1 => n18951, A2 => n18126, B1 => n18945, B2 => 
                           n17706, ZN => n6421);
   U3995 : OAI221_X1 port map( B1 => n3592, B2 => n18963, C1 => n18957, C2 => 
                           n2462, A => n6355, ZN => n6353);
   U3996 : AOI22_X1 port map( A1 => n18951, A2 => n18127, B1 => n18945, B2 => 
                           n17707, ZN => n6355);
   U3997 : OAI221_X1 port map( B1 => n3591, B2 => n18963, C1 => n18957, C2 => 
                           n2461, A => n6289, ZN => n6287);
   U3998 : AOI22_X1 port map( A1 => n18951, A2 => n18128, B1 => n18945, B2 => 
                           n17708, ZN => n6289);
   U3999 : OAI221_X1 port map( B1 => n3590, B2 => n18963, C1 => n18957, C2 => 
                           n2460, A => n6223, ZN => n6221);
   U4000 : AOI22_X1 port map( A1 => n18951, A2 => n18129, B1 => n18945, B2 => 
                           n17709, ZN => n6223);
   U4001 : OAI221_X1 port map( B1 => n3589, B2 => n18964, C1 => n18958, C2 => 
                           n2459, A => n6157, ZN => n6155);
   U4002 : AOI22_X1 port map( A1 => n18952, A2 => n18130, B1 => n18946, B2 => 
                           n17710, ZN => n6157);
   U4003 : OAI221_X1 port map( B1 => n3588, B2 => n18964, C1 => n18958, C2 => 
                           n2458, A => n6091, ZN => n6089);
   U4004 : AOI22_X1 port map( A1 => n18952, A2 => n18131, B1 => n18946, B2 => 
                           n17711, ZN => n6091);
   U4005 : OAI221_X1 port map( B1 => n3587, B2 => n18964, C1 => n18958, C2 => 
                           n2457, A => n6023, ZN => n6021);
   U4006 : AOI22_X1 port map( A1 => n18952, A2 => n18132, B1 => n18946, B2 => 
                           n17712, ZN => n6023);
   U4007 : OAI221_X1 port map( B1 => n3586, B2 => n18964, C1 => n18958, C2 => 
                           n2456, A => n5955, ZN => n5953);
   U4008 : AOI22_X1 port map( A1 => n18952, A2 => n18133, B1 => n18946, B2 => 
                           n17713, ZN => n5955);
   U4009 : OAI221_X1 port map( B1 => n3585, B2 => n18964, C1 => n18958, C2 => 
                           n2455, A => n5888, ZN => n5886);
   U4010 : AOI22_X1 port map( A1 => n18952, A2 => n18134, B1 => n18946, B2 => 
                           n17714, ZN => n5888);
   U4011 : OAI221_X1 port map( B1 => n3584, B2 => n18964, C1 => n18958, C2 => 
                           n2454, A => n5821, ZN => n5819);
   U4012 : AOI22_X1 port map( A1 => n18952, A2 => n18135, B1 => n18946, B2 => 
                           n17715, ZN => n5821);
   U4013 : OAI221_X1 port map( B1 => n3583, B2 => n18964, C1 => n18958, C2 => 
                           n2453, A => n5749, ZN => n5747);
   U4014 : AOI22_X1 port map( A1 => n18952, A2 => n18136, B1 => n18946, B2 => 
                           n17716, ZN => n5749);
   U4015 : OAI221_X1 port map( B1 => n3582, B2 => n18964, C1 => n18958, C2 => 
                           n2452, A => n5679, ZN => n5677);
   U4016 : AOI22_X1 port map( A1 => n18952, A2 => n18137, B1 => n18946, B2 => 
                           n17717, ZN => n5679);
   U4017 : OAI221_X1 port map( B1 => n3581, B2 => n18964, C1 => n18958, C2 => 
                           n2451, A => n5611, ZN => n5609);
   U4018 : AOI22_X1 port map( A1 => n18952, A2 => n18138, B1 => n18946, B2 => 
                           n17718, ZN => n5611);
   U4019 : OAI221_X1 port map( B1 => n3580, B2 => n18964, C1 => n18958, C2 => 
                           n2450, A => n5542, ZN => n5540);
   U4020 : AOI22_X1 port map( A1 => n18952, A2 => n18139, B1 => n18946, B2 => 
                           n17719, ZN => n5542);
   U4021 : OAI221_X1 port map( B1 => n3579, B2 => n18964, C1 => n18958, C2 => 
                           n2449, A => n5473, ZN => n5471);
   U4022 : AOI22_X1 port map( A1 => n18952, A2 => n18140, B1 => n18946, B2 => 
                           n17720, ZN => n5473);
   U4023 : OAI221_X1 port map( B1 => n3578, B2 => n18964, C1 => n18958, C2 => 
                           n2448, A => n5405, ZN => n5403);
   U4024 : AOI22_X1 port map( A1 => n18952, A2 => n18141, B1 => n18946, B2 => 
                           n17721, ZN => n5405);
   U4025 : OAI221_X1 port map( B1 => n3637, B2 => n18960, C1 => n18954, C2 => 
                           n2763, A => n11703, ZN => n11697);
   U4026 : AOI22_X1 port map( A1 => n18948, A2 => n11704, B1 => n18942, B2 => 
                           n11605, ZN => n11703);
   U4027 : OAI221_X1 port map( B1 => n3636, B2 => n18960, C1 => n18954, C2 => 
                           n2762, A => n11549, ZN => n11547);
   U4028 : AOI22_X1 port map( A1 => n18948, A2 => n11550, B1 => n18942, B2 => 
                           n11506, ZN => n11549);
   U4029 : OAI221_X1 port map( B1 => n3635, B2 => n18960, C1 => n18954, C2 => 
                           n2761, A => n11481, ZN => n11479);
   U4030 : AOI22_X1 port map( A1 => n18948, A2 => n11482, B1 => n18942, B2 => 
                           n11439, ZN => n11481);
   U4031 : OAI221_X1 port map( B1 => n3634, B2 => n18960, C1 => n18954, C2 => 
                           n2760, A => n11414, ZN => n11412);
   U4032 : AOI22_X1 port map( A1 => n18948, A2 => n11415, B1 => n18942, B2 => 
                           n11371, ZN => n11414);
   U4033 : OAI221_X1 port map( B1 => n3633, B2 => n18960, C1 => n18954, C2 => 
                           n2759, A => n11347, ZN => n11345);
   U4034 : AOI22_X1 port map( A1 => n18948, A2 => n18142, B1 => n18942, B2 => 
                           n17722, ZN => n11347);
   U4035 : OAI221_X1 port map( B1 => n3632, B2 => n18960, C1 => n18954, C2 => 
                           n2758, A => n11280, ZN => n11277);
   U4036 : AOI22_X1 port map( A1 => n18948, A2 => n18143, B1 => n18942, B2 => 
                           n17723, ZN => n11280);
   U4037 : OAI221_X1 port map( B1 => n3631, B2 => n18960, C1 => n18954, C2 => 
                           n2757, A => n11212, ZN => n11210);
   U4038 : AOI22_X1 port map( A1 => n18948, A2 => n18144, B1 => n18942, B2 => 
                           n17724, ZN => n11212);
   U4039 : OAI221_X1 port map( B1 => n3630, B2 => n18960, C1 => n18954, C2 => 
                           n2756, A => n11145, ZN => n11143);
   U4040 : AOI22_X1 port map( A1 => n18948, A2 => n18145, B1 => n18942, B2 => 
                           n17725, ZN => n11145);
   U4041 : OAI221_X1 port map( B1 => n3629, B2 => n18960, C1 => n18954, C2 => 
                           n2755, A => n11078, ZN => n11076);
   U4042 : AOI22_X1 port map( A1 => n18948, A2 => n18146, B1 => n18942, B2 => 
                           n17726, ZN => n11078);
   U4043 : OAI221_X1 port map( B1 => n3628, B2 => n18960, C1 => n18954, C2 => 
                           n2754, A => n11010, ZN => n11008);
   U4044 : AOI22_X1 port map( A1 => n18948, A2 => n18147, B1 => n18942, B2 => 
                           n17727, ZN => n11010);
   U4045 : OAI221_X1 port map( B1 => n3627, B2 => n18960, C1 => n18954, C2 => 
                           n2753, A => n10943, ZN => n10941);
   U4046 : AOI22_X1 port map( A1 => n18948, A2 => n18148, B1 => n18942, B2 => 
                           n17728, ZN => n10943);
   U4047 : OAI221_X1 port map( B1 => n3626, B2 => n18960, C1 => n18954, C2 => 
                           n2752, A => n10876, ZN => n10874);
   U4048 : AOI22_X1 port map( A1 => n18948, A2 => n18149, B1 => n18942, B2 => 
                           n17729, ZN => n10876);
   U4049 : OAI221_X1 port map( B1 => n3625, B2 => n18961, C1 => n18955, C2 => 
                           n2751, A => n10809, ZN => n10807);
   U4050 : AOI22_X1 port map( A1 => n18949, A2 => n18150, B1 => n18943, B2 => 
                           n17730, ZN => n10809);
   U4051 : OAI221_X1 port map( B1 => n3624, B2 => n18961, C1 => n18955, C2 => 
                           n2750, A => n10741, ZN => n10739);
   U4052 : AOI22_X1 port map( A1 => n18949, A2 => n18151, B1 => n18943, B2 => 
                           n17731, ZN => n10741);
   U4053 : OAI221_X1 port map( B1 => n3623, B2 => n18961, C1 => n18955, C2 => 
                           n2749, A => n10674, ZN => n10672);
   U4054 : AOI22_X1 port map( A1 => n18949, A2 => n18152, B1 => n18943, B2 => 
                           n17732, ZN => n10674);
   U4055 : OAI221_X1 port map( B1 => n3622, B2 => n18961, C1 => n18955, C2 => 
                           n2748, A => n10607, ZN => n10605);
   U4056 : AOI22_X1 port map( A1 => n18949, A2 => n18153, B1 => n18943, B2 => 
                           n17733, ZN => n10607);
   U4057 : OAI221_X1 port map( B1 => n3621, B2 => n18961, C1 => n18955, C2 => 
                           n2747, A => n10540, ZN => n10538);
   U4058 : AOI22_X1 port map( A1 => n18949, A2 => n18154, B1 => n18943, B2 => 
                           n17734, ZN => n10540);
   U4059 : OAI221_X1 port map( B1 => n3620, B2 => n18961, C1 => n18955, C2 => 
                           n2746, A => n10472, ZN => n10470);
   U4060 : AOI22_X1 port map( A1 => n18949, A2 => n18155, B1 => n18943, B2 => 
                           n17735, ZN => n10472);
   U4061 : OAI221_X1 port map( B1 => n3619, B2 => n18961, C1 => n18955, C2 => 
                           n2745, A => n10405, ZN => n10403);
   U4062 : AOI22_X1 port map( A1 => n18949, A2 => n18156, B1 => n18943, B2 => 
                           n17736, ZN => n10405);
   U4063 : OAI221_X1 port map( B1 => n3618, B2 => n18961, C1 => n18955, C2 => 
                           n2744, A => n10338, ZN => n10336);
   U4064 : AOI22_X1 port map( A1 => n18949, A2 => n18157, B1 => n18943, B2 => 
                           n17737, ZN => n10338);
   U4065 : OAI221_X1 port map( B1 => n3617, B2 => n18961, C1 => n18955, C2 => 
                           n2743, A => n10270, ZN => n10268);
   U4066 : AOI22_X1 port map( A1 => n18949, A2 => n18158, B1 => n18943, B2 => 
                           n17738, ZN => n10270);
   U4067 : OAI221_X1 port map( B1 => n3616, B2 => n18961, C1 => n18955, C2 => 
                           n2742, A => n10203, ZN => n10201);
   U4068 : AOI22_X1 port map( A1 => n18949, A2 => n18159, B1 => n18943, B2 => 
                           n17739, ZN => n10203);
   U4069 : OAI221_X1 port map( B1 => n3615, B2 => n18961, C1 => n18955, C2 => 
                           n2741, A => n10136, ZN => n10134);
   U4070 : AOI22_X1 port map( A1 => n18949, A2 => n18160, B1 => n18943, B2 => 
                           n17740, ZN => n10136);
   U4071 : OAI221_X1 port map( B1 => n3614, B2 => n18961, C1 => n18955, C2 => 
                           n2740, A => n10069, ZN => n10067);
   U4072 : AOI22_X1 port map( A1 => n18949, A2 => n18161, B1 => n18943, B2 => 
                           n17741, ZN => n10069);
   U4073 : OAI221_X1 port map( B1 => n3613, B2 => n18962, C1 => n18956, C2 => 
                           n2739, A => n10001, ZN => n9999);
   U4074 : AOI22_X1 port map( A1 => n18950, A2 => n18162, B1 => n18944, B2 => 
                           n17742, ZN => n10001);
   U4075 : OAI221_X1 port map( B1 => n3612, B2 => n18962, C1 => n18956, C2 => 
                           n2738, A => n9934, ZN => n9932);
   U4076 : AOI22_X1 port map( A1 => n18950, A2 => n18163, B1 => n18944, B2 => 
                           n17743, ZN => n9934);
   U4077 : OAI221_X1 port map( B1 => n3611, B2 => n18962, C1 => n18956, C2 => 
                           n2737, A => n9867, ZN => n9865);
   U4078 : AOI22_X1 port map( A1 => n18950, A2 => n18164, B1 => n18944, B2 => 
                           n17744, ZN => n9867);
   U4079 : OAI221_X1 port map( B1 => n3610, B2 => n18962, C1 => n18956, C2 => 
                           n2736, A => n9800, ZN => n9798);
   U4080 : AOI22_X1 port map( A1 => n18950, A2 => n18165, B1 => n18944, B2 => 
                           n17745, ZN => n9800);
   U4081 : OAI221_X1 port map( B1 => n3609, B2 => n18962, C1 => n18956, C2 => 
                           n2735, A => n9732, ZN => n9730);
   U4082 : AOI22_X1 port map( A1 => n18950, A2 => n18166, B1 => n18944, B2 => 
                           n17746, ZN => n9732);
   U4083 : OAI221_X1 port map( B1 => n3608, B2 => n18962, C1 => n18956, C2 => 
                           n2734, A => n9665, ZN => n9663);
   U4084 : AOI22_X1 port map( A1 => n18950, A2 => n18167, B1 => n18944, B2 => 
                           n17747, ZN => n9665);
   U4085 : OAI221_X1 port map( B1 => n3607, B2 => n18962, C1 => n18956, C2 => 
                           n2733, A => n9598, ZN => n9596);
   U4086 : AOI22_X1 port map( A1 => n18950, A2 => n18168, B1 => n18944, B2 => 
                           n17748, ZN => n9598);
   U4087 : OAI221_X1 port map( B1 => n3606, B2 => n18962, C1 => n18956, C2 => 
                           n2732, A => n9531, ZN => n9528);
   U4088 : AOI22_X1 port map( A1 => n18950, A2 => n18169, B1 => n18944, B2 => 
                           n17749, ZN => n9531);
   U4089 : OAI221_X1 port map( B1 => n3605, B2 => n18962, C1 => n18956, C2 => 
                           n2731, A => n9463, ZN => n9461);
   U4090 : AOI22_X1 port map( A1 => n18950, A2 => n18170, B1 => n18944, B2 => 
                           n17750, ZN => n9463);
   U4091 : OAI221_X1 port map( B1 => n3604, B2 => n18962, C1 => n18956, C2 => 
                           n2730, A => n9396, ZN => n9394);
   U4092 : AOI22_X1 port map( A1 => n18950, A2 => n18171, B1 => n18944, B2 => 
                           n17751, ZN => n9396);
   U4093 : OAI221_X1 port map( B1 => n3603, B2 => n18962, C1 => n18956, C2 => 
                           n2729, A => n9329, ZN => n9327);
   U4094 : AOI22_X1 port map( A1 => n18950, A2 => n18172, B1 => n18944, B2 => 
                           n17752, ZN => n9329);
   U4095 : OAI221_X1 port map( B1 => n3602, B2 => n18962, C1 => n18956, C2 => 
                           n2728, A => n7021, ZN => n7019);
   U4096 : AOI22_X1 port map( A1 => n18950, A2 => n18173, B1 => n18944, B2 => 
                           n17753, ZN => n7021);
   U4097 : OAI221_X1 port map( B1 => n3601, B2 => n18963, C1 => n18957, C2 => 
                           n2727, A => n6955, ZN => n6953);
   U4098 : AOI22_X1 port map( A1 => n18951, A2 => n18174, B1 => n18945, B2 => 
                           n17754, ZN => n6955);
   U4099 : OAI221_X1 port map( B1 => n3600, B2 => n18963, C1 => n18957, C2 => 
                           n2726, A => n6888, ZN => n6886);
   U4100 : AOI22_X1 port map( A1 => n18951, A2 => n18175, B1 => n18945, B2 => 
                           n17755, ZN => n6888);
   U4101 : OAI221_X1 port map( B1 => n4204, B2 => n19029, C1 => n1899, C2 => 
                           n19023, A => n6816, ZN => n6812);
   U4102 : AOI22_X1 port map( A1 => n19017, A2 => registers_15_38_port, B1 => 
                           n19011, B2 => n6785, ZN => n6816);
   U4103 : OAI221_X1 port map( B1 => n19005, B2 => n6760, C1 => n2122, C2 => 
                           n18999, A => n6817, ZN => n6811);
   U4104 : AOI22_X1 port map( A1 => n18993, A2 => n6818, B1 => n18987, B2 => 
                           registers_14_38_port, ZN => n6817);
   U4105 : OAI22_X1 port map( A1 => n5260, A2 => n19163, B1 => n3509, B2 => 
                           n19157, ZN => n5317);
   U4106 : OAI22_X1 port map( A1 => n5259, A2 => n19163, B1 => n3508, B2 => 
                           n19157, ZN => n4512);
   U4107 : OAI22_X1 port map( A1 => n5258, A2 => n19163, B1 => n3507, B2 => 
                           n19157, ZN => n3292);
   U4108 : OAI22_X1 port map( A1 => n5257, A2 => n19163, B1 => n3506, B2 => 
                           n19157, ZN => n3118);
   U4109 : OAI22_X1 port map( A1 => n5260, A2 => n19362, B1 => n3509, B2 => 
                           n19356, ZN => n5297);
   U4110 : OAI22_X1 port map( A1 => n5259, A2 => n19362, B1 => n3508, B2 => 
                           n19356, ZN => n4108);
   U4111 : OAI22_X1 port map( A1 => n5258, A2 => n19362, B1 => n3507, B2 => 
                           n19356, ZN => n3252);
   U4112 : OAI22_X1 port map( A1 => n5257, A2 => n19362, B1 => n3506, B2 => 
                           n19356, ZN => n3001);
   U4113 : OAI22_X1 port map( A1 => n4520, A2 => n18929, B1 => n4723, B2 => 
                           n18923, ZN => n5339);
   U4114 : OAI22_X1 port map( A1 => n4519, A2 => n18929, B1 => n4722, B2 => 
                           n18923, ZN => n4854);
   U4115 : OAI22_X1 port map( A1 => n4518, A2 => n18929, B1 => n4721, B2 => 
                           n18923, ZN => n3572);
   U4116 : OAI22_X1 port map( A1 => n4517, A2 => n18929, B1 => n4720, B2 => 
                           n18923, ZN => n3194);
   U4117 : OAI22_X1 port map( A1 => n4520, A2 => n19085, B1 => n4451, B2 => 
                           n19079, ZN => n5320);
   U4118 : OAI22_X1 port map( A1 => n4519, A2 => n19085, B1 => n4450, B2 => 
                           n19079, ZN => n4515);
   U4119 : OAI22_X1 port map( A1 => n4518, A2 => n19085, B1 => n4449, B2 => 
                           n19079, ZN => n3297);
   U4120 : OAI22_X1 port map( A1 => n4517, A2 => n19085, B1 => n4448, B2 => 
                           n19079, ZN => n3136);
   U4121 : OAI22_X1 port map( A1 => n4657, A2 => n19109, B1 => n3776, B2 => 
                           n19103, ZN => n5319);
   U4122 : OAI22_X1 port map( A1 => n4657, A2 => n19308, B1 => n3776, B2 => 
                           n19302, ZN => n5299);
   U4123 : OAI22_X1 port map( A1 => n4520, A2 => n19284, B1 => n4451, B2 => 
                           n19278, ZN => n5302);
   U4124 : OAI22_X1 port map( A1 => n4656, A2 => n19109, B1 => n3775, B2 => 
                           n19103, ZN => n4514);
   U4125 : OAI22_X1 port map( A1 => n4656, A2 => n19308, B1 => n3775, B2 => 
                           n19302, ZN => n4174);
   U4126 : OAI22_X1 port map( A1 => n4519, A2 => n19284, B1 => n4450, B2 => 
                           n19278, ZN => n4177);
   U4127 : OAI22_X1 port map( A1 => n4655, A2 => n19109, B1 => n3774, B2 => 
                           n19103, ZN => n3296);
   U4128 : OAI22_X1 port map( A1 => n4655, A2 => n19308, B1 => n3774, B2 => 
                           n19302, ZN => n3256);
   U4129 : OAI22_X1 port map( A1 => n4518, A2 => n19284, B1 => n4449, B2 => 
                           n19278, ZN => n3262);
   U4130 : OAI22_X1 port map( A1 => n4654, A2 => n19109, B1 => n3773, B2 => 
                           n19103, ZN => n3131);
   U4131 : OAI22_X1 port map( A1 => n4654, A2 => n19308, B1 => n3773, B2 => 
                           n19302, ZN => n3014);
   U4132 : OAI22_X1 port map( A1 => n4517, A2 => n19284, B1 => n4448, B2 => 
                           n19278, ZN => n3021);
   U4133 : OAI22_X1 port map( A1 => n6033, A2 => n19158, B1 => n3569, B2 => 
                           n19152, ZN => n11650);
   U4134 : OAI22_X1 port map( A1 => n6033, A2 => n19357, B1 => n3569, B2 => 
                           n19351, ZN => n11609);
   U4135 : OAI22_X1 port map( A1 => n5968, A2 => n19158, B1 => n3568, B2 => 
                           n19152, ZN => n11530);
   U4136 : OAI22_X1 port map( A1 => n5968, A2 => n19357, B1 => n3568, B2 => 
                           n19351, ZN => n11510);
   U4137 : OAI22_X1 port map( A1 => n5966, A2 => n19158, B1 => n3567, B2 => 
                           n19152, ZN => n11463);
   U4138 : OAI22_X1 port map( A1 => n5966, A2 => n19357, B1 => n3567, B2 => 
                           n19351, ZN => n11443);
   U4139 : OAI22_X1 port map( A1 => n5901, A2 => n19158, B1 => n3566, B2 => 
                           n19152, ZN => n11396);
   U4140 : OAI22_X1 port map( A1 => n5901, A2 => n19357, B1 => n3566, B2 => 
                           n19351, ZN => n11375);
   U4141 : OAI22_X1 port map( A1 => n5835, A2 => n19158, B1 => n3565, B2 => 
                           n19152, ZN => n11328);
   U4142 : OAI22_X1 port map( A1 => n5835, A2 => n19357, B1 => n3565, B2 => 
                           n19351, ZN => n11308);
   U4143 : OAI22_X1 port map( A1 => n5769, A2 => n19158, B1 => n3564, B2 => 
                           n19152, ZN => n11261);
   U4144 : OAI22_X1 port map( A1 => n5769, A2 => n19357, B1 => n3564, B2 => 
                           n19351, ZN => n11241);
   U4145 : OAI22_X1 port map( A1 => n5767, A2 => n19158, B1 => n3563, B2 => 
                           n19152, ZN => n11194);
   U4146 : OAI22_X1 port map( A1 => n5767, A2 => n19357, B1 => n3563, B2 => 
                           n19351, ZN => n11174);
   U4147 : OAI22_X1 port map( A1 => n5766, A2 => n19158, B1 => n3562, B2 => 
                           n19152, ZN => n11127);
   U4148 : OAI22_X1 port map( A1 => n5766, A2 => n19357, B1 => n3562, B2 => 
                           n19351, ZN => n11106);
   U4149 : OAI22_X1 port map( A1 => n5765, A2 => n19158, B1 => n3561, B2 => 
                           n19152, ZN => n11059);
   U4150 : OAI22_X1 port map( A1 => n5765, A2 => n19357, B1 => n3561, B2 => 
                           n19351, ZN => n11039);
   U4151 : OAI22_X1 port map( A1 => n5764, A2 => n19158, B1 => n3560, B2 => 
                           n19152, ZN => n10992);
   U4152 : OAI22_X1 port map( A1 => n5764, A2 => n19357, B1 => n3560, B2 => 
                           n19351, ZN => n10972);
   U4153 : OAI22_X1 port map( A1 => n5763, A2 => n19158, B1 => n3559, B2 => 
                           n19152, ZN => n10925);
   U4154 : OAI22_X1 port map( A1 => n5763, A2 => n19357, B1 => n3559, B2 => 
                           n19351, ZN => n10904);
   U4155 : OAI22_X1 port map( A1 => n5698, A2 => n19158, B1 => n3558, B2 => 
                           n19152, ZN => n10858);
   U4156 : OAI22_X1 port map( A1 => n5698, A2 => n19357, B1 => n3558, B2 => 
                           n19351, ZN => n10837);
   U4157 : OAI22_X1 port map( A1 => n5696, A2 => n19159, B1 => n3557, B2 => 
                           n19153, ZN => n10790);
   U4158 : OAI22_X1 port map( A1 => n5696, A2 => n19358, B1 => n3557, B2 => 
                           n19352, ZN => n10770);
   U4159 : OAI22_X1 port map( A1 => n5695, A2 => n19159, B1 => n3556, B2 => 
                           n19153, ZN => n10723);
   U4160 : OAI22_X1 port map( A1 => n5695, A2 => n19358, B1 => n3556, B2 => 
                           n19352, ZN => n10703);
   U4161 : OAI22_X1 port map( A1 => n5694, A2 => n19159, B1 => n3555, B2 => 
                           n19153, ZN => n10656);
   U4162 : OAI22_X1 port map( A1 => n5694, A2 => n19358, B1 => n3555, B2 => 
                           n19352, ZN => n10635);
   U4163 : OAI22_X1 port map( A1 => n5629, A2 => n19159, B1 => n3554, B2 => 
                           n19153, ZN => n10588);
   U4164 : OAI22_X1 port map( A1 => n5629, A2 => n19358, B1 => n3554, B2 => 
                           n19352, ZN => n10568);
   U4165 : OAI22_X1 port map( A1 => n5627, A2 => n19159, B1 => n3553, B2 => 
                           n19153, ZN => n10521);
   U4166 : OAI22_X1 port map( A1 => n5627, A2 => n19358, B1 => n3553, B2 => 
                           n19352, ZN => n10501);
   U4167 : OAI22_X1 port map( A1 => n5562, A2 => n19159, B1 => n3552, B2 => 
                           n19153, ZN => n10454);
   U4168 : OAI22_X1 port map( A1 => n5562, A2 => n19358, B1 => n3552, B2 => 
                           n19352, ZN => n10434);
   U4169 : OAI22_X1 port map( A1 => n5560, A2 => n19159, B1 => n3551, B2 => 
                           n19153, ZN => n10387);
   U4170 : OAI22_X1 port map( A1 => n5560, A2 => n19358, B1 => n3551, B2 => 
                           n19352, ZN => n10366);
   U4171 : OAI22_X1 port map( A1 => n5559, A2 => n19159, B1 => n3550, B2 => 
                           n19153, ZN => n10319);
   U4172 : OAI22_X1 port map( A1 => n5559, A2 => n19358, B1 => n3550, B2 => 
                           n19352, ZN => n10299);
   U4173 : OAI22_X1 port map( A1 => n5494, A2 => n19159, B1 => n3549, B2 => 
                           n19153, ZN => n10252);
   U4174 : OAI22_X1 port map( A1 => n5494, A2 => n19358, B1 => n3549, B2 => 
                           n19352, ZN => n10232);
   U4175 : OAI22_X1 port map( A1 => n5492, A2 => n19159, B1 => n3548, B2 => 
                           n19153, ZN => n10185);
   U4176 : OAI22_X1 port map( A1 => n5492, A2 => n19358, B1 => n3548, B2 => 
                           n19352, ZN => n10164);
   U4177 : OAI22_X1 port map( A1 => n5491, A2 => n19159, B1 => n3547, B2 => 
                           n19153, ZN => n10118);
   U4178 : OAI22_X1 port map( A1 => n5491, A2 => n19358, B1 => n3547, B2 => 
                           n19352, ZN => n10097);
   U4179 : OAI22_X1 port map( A1 => n5426, A2 => n19159, B1 => n3546, B2 => 
                           n19153, ZN => n10050);
   U4180 : OAI22_X1 port map( A1 => n5426, A2 => n19358, B1 => n3546, B2 => 
                           n19352, ZN => n10030);
   U4181 : OAI22_X1 port map( A1 => n5424, A2 => n19160, B1 => n3545, B2 => 
                           n19154, ZN => n9983);
   U4182 : OAI22_X1 port map( A1 => n5424, A2 => n19359, B1 => n3545, B2 => 
                           n19353, ZN => n9963);
   U4183 : OAI22_X1 port map( A1 => n5359, A2 => n19160, B1 => n3544, B2 => 
                           n19154, ZN => n9916);
   U4184 : OAI22_X1 port map( A1 => n5359, A2 => n19359, B1 => n3544, B2 => 
                           n19353, ZN => n9895);
   U4185 : OAI22_X1 port map( A1 => n5357, A2 => n19160, B1 => n3543, B2 => 
                           n19154, ZN => n9849);
   U4186 : OAI22_X1 port map( A1 => n5357, A2 => n19359, B1 => n3543, B2 => 
                           n19353, ZN => n9828);
   U4187 : OAI22_X1 port map( A1 => n5356, A2 => n19160, B1 => n3542, B2 => 
                           n19154, ZN => n9781);
   U4188 : OAI22_X1 port map( A1 => n5356, A2 => n19359, B1 => n3542, B2 => 
                           n19353, ZN => n9761);
   U4189 : OAI22_X1 port map( A1 => n5355, A2 => n19160, B1 => n3541, B2 => 
                           n19154, ZN => n9714);
   U4190 : OAI22_X1 port map( A1 => n5355, A2 => n19359, B1 => n3541, B2 => 
                           n19353, ZN => n9694);
   U4191 : OAI22_X1 port map( A1 => n5291, A2 => n19160, B1 => n3540, B2 => 
                           n19154, ZN => n9647);
   U4192 : OAI22_X1 port map( A1 => n5291, A2 => n19359, B1 => n3540, B2 => 
                           n19353, ZN => n9626);
   U4193 : OAI22_X1 port map( A1 => n5290, A2 => n19160, B1 => n3539, B2 => 
                           n19154, ZN => n9579);
   U4194 : OAI22_X1 port map( A1 => n5290, A2 => n19359, B1 => n3539, B2 => 
                           n19353, ZN => n9559);
   U4195 : OAI22_X1 port map( A1 => n5289, A2 => n19160, B1 => n3538, B2 => 
                           n19154, ZN => n9512);
   U4196 : OAI22_X1 port map( A1 => n5289, A2 => n19359, B1 => n3538, B2 => 
                           n19353, ZN => n9492);
   U4197 : OAI22_X1 port map( A1 => n5288, A2 => n19160, B1 => n3537, B2 => 
                           n19154, ZN => n9445);
   U4198 : OAI22_X1 port map( A1 => n5288, A2 => n19359, B1 => n3537, B2 => 
                           n19353, ZN => n9425);
   U4199 : OAI22_X1 port map( A1 => n5287, A2 => n19160, B1 => n3536, B2 => 
                           n19154, ZN => n9378);
   U4200 : OAI22_X1 port map( A1 => n5287, A2 => n19359, B1 => n3536, B2 => 
                           n19353, ZN => n9357);
   U4201 : OAI22_X1 port map( A1 => n5286, A2 => n19160, B1 => n3535, B2 => 
                           n19154, ZN => n9310);
   U4202 : OAI22_X1 port map( A1 => n5286, A2 => n19359, B1 => n3535, B2 => 
                           n19353, ZN => n9290);
   U4203 : OAI22_X1 port map( A1 => n5285, A2 => n19160, B1 => n3534, B2 => 
                           n19154, ZN => n7003);
   U4204 : OAI22_X1 port map( A1 => n5285, A2 => n19359, B1 => n3534, B2 => 
                           n19353, ZN => n6983);
   U4205 : OAI22_X1 port map( A1 => n5284, A2 => n19161, B1 => n3533, B2 => 
                           n19155, ZN => n6936);
   U4206 : OAI22_X1 port map( A1 => n5284, A2 => n19360, B1 => n3533, B2 => 
                           n19354, ZN => n6916);
   U4207 : OAI22_X1 port map( A1 => n5283, A2 => n19161, B1 => n3532, B2 => 
                           n19155, ZN => n6870);
   U4208 : OAI22_X1 port map( A1 => n5283, A2 => n19360, B1 => n3532, B2 => 
                           n19354, ZN => n6849);
   U4209 : OAI22_X1 port map( A1 => n5282, A2 => n19161, B1 => n3531, B2 => 
                           n19155, ZN => n6803);
   U4210 : OAI22_X1 port map( A1 => n5282, A2 => n19360, B1 => n3531, B2 => 
                           n19354, ZN => n6782);
   U4211 : OAI22_X1 port map( A1 => n5281, A2 => n19161, B1 => n3530, B2 => 
                           n19155, ZN => n6735);
   U4212 : OAI22_X1 port map( A1 => n5281, A2 => n19360, B1 => n3530, B2 => 
                           n19354, ZN => n6715);
   U4213 : OAI22_X1 port map( A1 => n5280, A2 => n19161, B1 => n3529, B2 => 
                           n19155, ZN => n6668);
   U4214 : OAI22_X1 port map( A1 => n5280, A2 => n19360, B1 => n3529, B2 => 
                           n19354, ZN => n6648);
   U4215 : OAI22_X1 port map( A1 => n5279, A2 => n19161, B1 => n3528, B2 => 
                           n19155, ZN => n6601);
   U4216 : OAI22_X1 port map( A1 => n5279, A2 => n19360, B1 => n3528, B2 => 
                           n19354, ZN => n6581);
   U4217 : OAI22_X1 port map( A1 => n5278, A2 => n19161, B1 => n3527, B2 => 
                           n19155, ZN => n6535);
   U4218 : OAI22_X1 port map( A1 => n5278, A2 => n19360, B1 => n3527, B2 => 
                           n19354, ZN => n6515);
   U4219 : OAI22_X1 port map( A1 => n5277, A2 => n19161, B1 => n3526, B2 => 
                           n19155, ZN => n6469);
   U4220 : OAI22_X1 port map( A1 => n5277, A2 => n19360, B1 => n3526, B2 => 
                           n19354, ZN => n6449);
   U4221 : OAI22_X1 port map( A1 => n5276, A2 => n19161, B1 => n3525, B2 => 
                           n19155, ZN => n6403);
   U4222 : OAI22_X1 port map( A1 => n5276, A2 => n19360, B1 => n3525, B2 => 
                           n19354, ZN => n6383);
   U4223 : OAI22_X1 port map( A1 => n5275, A2 => n19161, B1 => n3524, B2 => 
                           n19155, ZN => n6337);
   U4224 : OAI22_X1 port map( A1 => n5275, A2 => n19360, B1 => n3524, B2 => 
                           n19354, ZN => n6317);
   U4225 : OAI22_X1 port map( A1 => n5274, A2 => n19161, B1 => n3523, B2 => 
                           n19155, ZN => n6271);
   U4226 : OAI22_X1 port map( A1 => n5274, A2 => n19360, B1 => n3523, B2 => 
                           n19354, ZN => n6251);
   U4227 : OAI22_X1 port map( A1 => n5273, A2 => n19161, B1 => n3522, B2 => 
                           n19155, ZN => n6205);
   U4228 : OAI22_X1 port map( A1 => n5273, A2 => n19360, B1 => n3522, B2 => 
                           n19354, ZN => n6185);
   U4229 : OAI22_X1 port map( A1 => n5272, A2 => n19162, B1 => n3521, B2 => 
                           n19156, ZN => n6139);
   U4230 : OAI22_X1 port map( A1 => n5272, A2 => n19361, B1 => n3521, B2 => 
                           n19355, ZN => n6119);
   U4231 : OAI22_X1 port map( A1 => n5271, A2 => n19162, B1 => n3520, B2 => 
                           n19156, ZN => n6073);
   U4232 : OAI22_X1 port map( A1 => n5271, A2 => n19361, B1 => n3520, B2 => 
                           n19355, ZN => n6053);
   U4233 : OAI22_X1 port map( A1 => n5270, A2 => n19162, B1 => n3519, B2 => 
                           n19156, ZN => n6005);
   U4234 : OAI22_X1 port map( A1 => n5270, A2 => n19361, B1 => n3519, B2 => 
                           n19355, ZN => n5985);
   U4235 : OAI22_X1 port map( A1 => n5269, A2 => n19162, B1 => n3518, B2 => 
                           n19156, ZN => n5937);
   U4236 : OAI22_X1 port map( A1 => n5269, A2 => n19361, B1 => n3518, B2 => 
                           n19355, ZN => n5917);
   U4237 : OAI22_X1 port map( A1 => n5268, A2 => n19162, B1 => n3517, B2 => 
                           n19156, ZN => n5870);
   U4238 : OAI22_X1 port map( A1 => n5268, A2 => n19361, B1 => n3517, B2 => 
                           n19355, ZN => n5850);
   U4239 : OAI22_X1 port map( A1 => n5267, A2 => n19162, B1 => n3516, B2 => 
                           n19156, ZN => n5803);
   U4240 : OAI22_X1 port map( A1 => n5267, A2 => n19361, B1 => n3516, B2 => 
                           n19355, ZN => n5783);
   U4241 : OAI22_X1 port map( A1 => n5266, A2 => n19162, B1 => n3515, B2 => 
                           n19156, ZN => n5731);
   U4242 : OAI22_X1 port map( A1 => n5266, A2 => n19361, B1 => n3515, B2 => 
                           n19355, ZN => n5711);
   U4243 : OAI22_X1 port map( A1 => n5265, A2 => n19162, B1 => n3514, B2 => 
                           n19156, ZN => n5661);
   U4244 : OAI22_X1 port map( A1 => n5265, A2 => n19361, B1 => n3514, B2 => 
                           n19355, ZN => n5641);
   U4245 : OAI22_X1 port map( A1 => n5264, A2 => n19162, B1 => n3513, B2 => 
                           n19156, ZN => n5593);
   U4246 : OAI22_X1 port map( A1 => n5264, A2 => n19361, B1 => n3513, B2 => 
                           n19355, ZN => n5573);
   U4247 : OAI22_X1 port map( A1 => n5263, A2 => n19162, B1 => n3512, B2 => 
                           n19156, ZN => n5524);
   U4248 : OAI22_X1 port map( A1 => n5263, A2 => n19361, B1 => n3512, B2 => 
                           n19355, ZN => n5504);
   U4249 : OAI22_X1 port map( A1 => n5262, A2 => n19162, B1 => n3511, B2 => 
                           n19156, ZN => n5455);
   U4250 : OAI22_X1 port map( A1 => n5262, A2 => n19361, B1 => n3511, B2 => 
                           n19355, ZN => n5435);
   U4251 : OAI22_X1 port map( A1 => n5261, A2 => n19162, B1 => n3510, B2 => 
                           n19156, ZN => n5387);
   U4252 : OAI22_X1 port map( A1 => n5261, A2 => n19361, B1 => n3510, B2 => 
                           n19355, ZN => n5367);
   U4253 : OAI22_X1 port map( A1 => n4927, A2 => n18977, B1 => n4993, B2 => 
                           n18971, ZN => n5334);
   U4254 : OAI22_X1 port map( A1 => n4926, A2 => n18977, B1 => n4992, B2 => 
                           n18971, ZN => n4785);
   U4255 : OAI22_X1 port map( A1 => n4925, A2 => n18977, B1 => n4991, B2 => 
                           n18971, ZN => n3503);
   U4256 : OAI22_X1 port map( A1 => n4924, A2 => n18977, B1 => n4990, B2 => 
                           n18971, ZN => n3168);
   U4257 : OAI22_X1 port map( A1 => n4717, A2 => n19104, B1 => n3836, B2 => 
                           n19098, ZN => n11657);
   U4258 : OAI22_X1 port map( A1 => n4717, A2 => n19303, B1 => n3836, B2 => 
                           n19297, ZN => n11615);
   U4259 : OAI22_X1 port map( A1 => n4716, A2 => n19104, B1 => n3835, B2 => 
                           n19098, ZN => n11532);
   U4260 : OAI22_X1 port map( A1 => n4716, A2 => n19303, B1 => n3835, B2 => 
                           n19297, ZN => n11512);
   U4261 : OAI22_X1 port map( A1 => n4715, A2 => n19104, B1 => n3834, B2 => 
                           n19098, ZN => n11465);
   U4262 : OAI22_X1 port map( A1 => n4715, A2 => n19303, B1 => n3834, B2 => 
                           n19297, ZN => n11445);
   U4263 : OAI22_X1 port map( A1 => n4714, A2 => n19104, B1 => n3833, B2 => 
                           n19098, ZN => n11398);
   U4264 : OAI22_X1 port map( A1 => n4714, A2 => n19303, B1 => n3833, B2 => 
                           n19297, ZN => n11377);
   U4265 : OAI22_X1 port map( A1 => n4713, A2 => n19104, B1 => n3832, B2 => 
                           n19098, ZN => n11330);
   U4266 : OAI22_X1 port map( A1 => n4713, A2 => n19303, B1 => n3832, B2 => 
                           n19297, ZN => n11310);
   U4267 : OAI22_X1 port map( A1 => n4712, A2 => n19104, B1 => n3831, B2 => 
                           n19098, ZN => n11263);
   U4268 : OAI22_X1 port map( A1 => n4712, A2 => n19303, B1 => n3831, B2 => 
                           n19297, ZN => n11243);
   U4269 : OAI22_X1 port map( A1 => n4711, A2 => n19104, B1 => n3830, B2 => 
                           n19098, ZN => n11196);
   U4270 : OAI22_X1 port map( A1 => n4711, A2 => n19303, B1 => n3830, B2 => 
                           n19297, ZN => n11176);
   U4271 : OAI22_X1 port map( A1 => n4710, A2 => n19104, B1 => n3829, B2 => 
                           n19098, ZN => n11129);
   U4272 : OAI22_X1 port map( A1 => n4710, A2 => n19303, B1 => n3829, B2 => 
                           n19297, ZN => n11108);
   U4273 : OAI22_X1 port map( A1 => n4709, A2 => n19104, B1 => n3828, B2 => 
                           n19098, ZN => n11061);
   U4274 : OAI22_X1 port map( A1 => n4709, A2 => n19303, B1 => n3828, B2 => 
                           n19297, ZN => n11041);
   U4275 : OAI22_X1 port map( A1 => n4708, A2 => n19104, B1 => n3827, B2 => 
                           n19098, ZN => n10994);
   U4276 : OAI22_X1 port map( A1 => n4708, A2 => n19303, B1 => n3827, B2 => 
                           n19297, ZN => n10974);
   U4277 : OAI22_X1 port map( A1 => n4707, A2 => n19104, B1 => n3826, B2 => 
                           n19098, ZN => n10927);
   U4278 : OAI22_X1 port map( A1 => n4707, A2 => n19303, B1 => n3826, B2 => 
                           n19297, ZN => n10906);
   U4279 : OAI22_X1 port map( A1 => n4706, A2 => n19104, B1 => n3825, B2 => 
                           n19098, ZN => n10860);
   U4280 : OAI22_X1 port map( A1 => n4706, A2 => n19303, B1 => n3825, B2 => 
                           n19297, ZN => n10839);
   U4281 : OAI22_X1 port map( A1 => n4705, A2 => n19105, B1 => n3824, B2 => 
                           n19099, ZN => n10792);
   U4282 : OAI22_X1 port map( A1 => n4705, A2 => n19304, B1 => n3824, B2 => 
                           n19298, ZN => n10772);
   U4283 : OAI22_X1 port map( A1 => n4704, A2 => n19105, B1 => n3823, B2 => 
                           n19099, ZN => n10725);
   U4284 : OAI22_X1 port map( A1 => n4704, A2 => n19304, B1 => n3823, B2 => 
                           n19298, ZN => n10705);
   U4285 : OAI22_X1 port map( A1 => n4703, A2 => n19105, B1 => n3822, B2 => 
                           n19099, ZN => n10658);
   U4286 : OAI22_X1 port map( A1 => n4703, A2 => n19304, B1 => n3822, B2 => 
                           n19298, ZN => n10637);
   U4287 : OAI22_X1 port map( A1 => n4702, A2 => n19105, B1 => n3821, B2 => 
                           n19099, ZN => n10591);
   U4288 : OAI22_X1 port map( A1 => n4702, A2 => n19304, B1 => n3821, B2 => 
                           n19298, ZN => n10570);
   U4289 : OAI22_X1 port map( A1 => n4701, A2 => n19105, B1 => n3820, B2 => 
                           n19099, ZN => n10523);
   U4290 : OAI22_X1 port map( A1 => n4701, A2 => n19304, B1 => n3820, B2 => 
                           n19298, ZN => n10503);
   U4291 : OAI22_X1 port map( A1 => n4700, A2 => n19105, B1 => n3819, B2 => 
                           n19099, ZN => n10456);
   U4292 : OAI22_X1 port map( A1 => n4700, A2 => n19304, B1 => n3819, B2 => 
                           n19298, ZN => n10436);
   U4293 : OAI22_X1 port map( A1 => n4699, A2 => n19105, B1 => n3818, B2 => 
                           n19099, ZN => n10389);
   U4294 : OAI22_X1 port map( A1 => n4699, A2 => n19304, B1 => n3818, B2 => 
                           n19298, ZN => n10368);
   U4295 : OAI22_X1 port map( A1 => n4698, A2 => n19105, B1 => n3817, B2 => 
                           n19099, ZN => n10321);
   U4296 : OAI22_X1 port map( A1 => n4698, A2 => n19304, B1 => n3817, B2 => 
                           n19298, ZN => n10301);
   U4297 : OAI22_X1 port map( A1 => n4697, A2 => n19105, B1 => n3816, B2 => 
                           n19099, ZN => n10254);
   U4298 : OAI22_X1 port map( A1 => n4697, A2 => n19304, B1 => n3816, B2 => 
                           n19298, ZN => n10234);
   U4299 : OAI22_X1 port map( A1 => n4696, A2 => n19105, B1 => n3815, B2 => 
                           n19099, ZN => n10187);
   U4300 : OAI22_X1 port map( A1 => n4696, A2 => n19304, B1 => n3815, B2 => 
                           n19298, ZN => n10167);
   U4301 : OAI22_X1 port map( A1 => n4695, A2 => n19105, B1 => n3814, B2 => 
                           n19099, ZN => n10120);
   U4302 : OAI22_X1 port map( A1 => n4695, A2 => n19304, B1 => n3814, B2 => 
                           n19298, ZN => n10099);
   U4303 : OAI22_X1 port map( A1 => n4694, A2 => n19105, B1 => n3813, B2 => 
                           n19099, ZN => n10052);
   U4304 : OAI22_X1 port map( A1 => n4694, A2 => n19304, B1 => n3813, B2 => 
                           n19298, ZN => n10032);
   U4305 : OAI22_X1 port map( A1 => n4693, A2 => n19106, B1 => n3812, B2 => 
                           n19100, ZN => n9985);
   U4306 : OAI22_X1 port map( A1 => n4693, A2 => n19305, B1 => n3812, B2 => 
                           n19299, ZN => n9965);
   U4307 : OAI22_X1 port map( A1 => n4692, A2 => n19106, B1 => n3811, B2 => 
                           n19100, ZN => n9918);
   U4308 : OAI22_X1 port map( A1 => n4692, A2 => n19305, B1 => n3811, B2 => 
                           n19299, ZN => n9897);
   U4309 : OAI22_X1 port map( A1 => n4691, A2 => n19106, B1 => n3810, B2 => 
                           n19100, ZN => n9851);
   U4310 : OAI22_X1 port map( A1 => n4691, A2 => n19305, B1 => n3810, B2 => 
                           n19299, ZN => n9830);
   U4311 : OAI22_X1 port map( A1 => n4690, A2 => n19106, B1 => n3809, B2 => 
                           n19100, ZN => n9783);
   U4312 : OAI22_X1 port map( A1 => n4690, A2 => n19305, B1 => n3809, B2 => 
                           n19299, ZN => n9763);
   U4313 : OAI22_X1 port map( A1 => n4689, A2 => n19106, B1 => n3808, B2 => 
                           n19100, ZN => n9716);
   U4314 : OAI22_X1 port map( A1 => n4689, A2 => n19305, B1 => n3808, B2 => 
                           n19299, ZN => n9696);
   U4315 : OAI22_X1 port map( A1 => n4688, A2 => n19106, B1 => n3807, B2 => 
                           n19100, ZN => n9649);
   U4316 : OAI22_X1 port map( A1 => n4688, A2 => n19305, B1 => n3807, B2 => 
                           n19299, ZN => n9628);
   U4317 : OAI22_X1 port map( A1 => n4687, A2 => n19106, B1 => n3806, B2 => 
                           n19100, ZN => n9581);
   U4318 : OAI22_X1 port map( A1 => n4687, A2 => n19305, B1 => n3806, B2 => 
                           n19299, ZN => n9561);
   U4319 : OAI22_X1 port map( A1 => n4686, A2 => n19106, B1 => n3805, B2 => 
                           n19100, ZN => n9514);
   U4320 : OAI22_X1 port map( A1 => n4686, A2 => n19305, B1 => n3805, B2 => 
                           n19299, ZN => n9494);
   U4321 : OAI22_X1 port map( A1 => n4685, A2 => n19106, B1 => n3804, B2 => 
                           n19100, ZN => n9447);
   U4322 : OAI22_X1 port map( A1 => n4685, A2 => n19305, B1 => n3804, B2 => 
                           n19299, ZN => n9427);
   U4323 : OAI22_X1 port map( A1 => n4684, A2 => n19106, B1 => n3803, B2 => 
                           n19100, ZN => n9380);
   U4324 : OAI22_X1 port map( A1 => n4684, A2 => n19305, B1 => n3803, B2 => 
                           n19299, ZN => n9359);
   U4325 : OAI22_X1 port map( A1 => n4683, A2 => n19106, B1 => n3802, B2 => 
                           n19100, ZN => n9312);
   U4326 : OAI22_X1 port map( A1 => n4683, A2 => n19305, B1 => n3802, B2 => 
                           n19299, ZN => n9292);
   U4327 : OAI22_X1 port map( A1 => n4682, A2 => n19106, B1 => n3801, B2 => 
                           n19100, ZN => n7005);
   U4328 : OAI22_X1 port map( A1 => n4682, A2 => n19305, B1 => n3801, B2 => 
                           n19299, ZN => n6985);
   U4329 : OAI22_X1 port map( A1 => n4681, A2 => n19107, B1 => n3800, B2 => 
                           n19101, ZN => n6938);
   U4330 : OAI22_X1 port map( A1 => n4681, A2 => n19306, B1 => n3800, B2 => 
                           n19300, ZN => n6918);
   U4331 : OAI22_X1 port map( A1 => n4680, A2 => n19107, B1 => n3799, B2 => 
                           n19101, ZN => n6872);
   U4332 : OAI22_X1 port map( A1 => n4680, A2 => n19306, B1 => n3799, B2 => 
                           n19300, ZN => n6851);
   U4333 : OAI22_X1 port map( A1 => n4679, A2 => n19107, B1 => n3798, B2 => 
                           n19101, ZN => n6805);
   U4334 : OAI22_X1 port map( A1 => n4679, A2 => n19306, B1 => n3798, B2 => 
                           n19300, ZN => n6784);
   U4335 : OAI22_X1 port map( A1 => n4678, A2 => n19107, B1 => n3797, B2 => 
                           n19101, ZN => n6737);
   U4336 : OAI22_X1 port map( A1 => n4678, A2 => n19306, B1 => n3797, B2 => 
                           n19300, ZN => n6717);
   U4337 : OAI22_X1 port map( A1 => n4677, A2 => n19107, B1 => n3796, B2 => 
                           n19101, ZN => n6670);
   U4338 : OAI22_X1 port map( A1 => n4677, A2 => n19306, B1 => n3796, B2 => 
                           n19300, ZN => n6650);
   U4339 : OAI22_X1 port map( A1 => n4676, A2 => n19107, B1 => n3795, B2 => 
                           n19101, ZN => n6603);
   U4340 : OAI22_X1 port map( A1 => n4676, A2 => n19306, B1 => n3795, B2 => 
                           n19300, ZN => n6583);
   U4341 : OAI22_X1 port map( A1 => n4675, A2 => n19107, B1 => n3794, B2 => 
                           n19101, ZN => n6537);
   U4342 : OAI22_X1 port map( A1 => n4675, A2 => n19306, B1 => n3794, B2 => 
                           n19300, ZN => n6517);
   U4343 : OAI22_X1 port map( A1 => n4674, A2 => n19107, B1 => n3793, B2 => 
                           n19101, ZN => n6471);
   U4344 : OAI22_X1 port map( A1 => n4674, A2 => n19306, B1 => n3793, B2 => 
                           n19300, ZN => n6451);
   U4345 : OAI22_X1 port map( A1 => n4673, A2 => n19107, B1 => n3792, B2 => 
                           n19101, ZN => n6405);
   U4346 : OAI22_X1 port map( A1 => n4673, A2 => n19306, B1 => n3792, B2 => 
                           n19300, ZN => n6385);
   U4347 : OAI22_X1 port map( A1 => n4672, A2 => n19107, B1 => n3791, B2 => 
                           n19101, ZN => n6339);
   U4348 : OAI22_X1 port map( A1 => n4672, A2 => n19306, B1 => n3791, B2 => 
                           n19300, ZN => n6319);
   U4349 : OAI22_X1 port map( A1 => n4671, A2 => n19107, B1 => n3790, B2 => 
                           n19101, ZN => n6273);
   U4350 : OAI22_X1 port map( A1 => n4671, A2 => n19306, B1 => n3790, B2 => 
                           n19300, ZN => n6253);
   U4351 : OAI22_X1 port map( A1 => n4670, A2 => n19107, B1 => n3789, B2 => 
                           n19101, ZN => n6207);
   U4352 : OAI22_X1 port map( A1 => n4670, A2 => n19306, B1 => n3789, B2 => 
                           n19300, ZN => n6187);
   U4353 : OAI22_X1 port map( A1 => n4669, A2 => n19108, B1 => n3788, B2 => 
                           n19102, ZN => n6141);
   U4354 : OAI22_X1 port map( A1 => n4669, A2 => n19307, B1 => n3788, B2 => 
                           n19301, ZN => n6121);
   U4355 : OAI22_X1 port map( A1 => n4668, A2 => n19108, B1 => n3787, B2 => 
                           n19102, ZN => n6075);
   U4356 : OAI22_X1 port map( A1 => n4668, A2 => n19307, B1 => n3787, B2 => 
                           n19301, ZN => n6055);
   U4357 : OAI22_X1 port map( A1 => n4667, A2 => n19108, B1 => n3786, B2 => 
                           n19102, ZN => n6007);
   U4358 : OAI22_X1 port map( A1 => n4667, A2 => n19307, B1 => n3786, B2 => 
                           n19301, ZN => n5987);
   U4359 : OAI22_X1 port map( A1 => n4666, A2 => n19108, B1 => n3785, B2 => 
                           n19102, ZN => n5939);
   U4360 : OAI22_X1 port map( A1 => n4666, A2 => n19307, B1 => n3785, B2 => 
                           n19301, ZN => n5919);
   U4361 : OAI22_X1 port map( A1 => n4665, A2 => n19108, B1 => n3784, B2 => 
                           n19102, ZN => n5872);
   U4362 : OAI22_X1 port map( A1 => n4665, A2 => n19307, B1 => n3784, B2 => 
                           n19301, ZN => n5852);
   U4363 : OAI22_X1 port map( A1 => n4664, A2 => n19108, B1 => n3783, B2 => 
                           n19102, ZN => n5805);
   U4364 : OAI22_X1 port map( A1 => n4664, A2 => n19307, B1 => n3783, B2 => 
                           n19301, ZN => n5785);
   U4365 : OAI22_X1 port map( A1 => n4663, A2 => n19108, B1 => n3782, B2 => 
                           n19102, ZN => n5733);
   U4366 : OAI22_X1 port map( A1 => n4663, A2 => n19307, B1 => n3782, B2 => 
                           n19301, ZN => n5713);
   U4367 : OAI22_X1 port map( A1 => n4662, A2 => n19108, B1 => n3781, B2 => 
                           n19102, ZN => n5663);
   U4368 : OAI22_X1 port map( A1 => n4662, A2 => n19307, B1 => n3781, B2 => 
                           n19301, ZN => n5643);
   U4369 : OAI22_X1 port map( A1 => n4661, A2 => n19108, B1 => n3780, B2 => 
                           n19102, ZN => n5595);
   U4370 : OAI22_X1 port map( A1 => n4661, A2 => n19307, B1 => n3780, B2 => 
                           n19301, ZN => n5575);
   U4371 : OAI22_X1 port map( A1 => n4660, A2 => n19108, B1 => n3779, B2 => 
                           n19102, ZN => n5526);
   U4372 : OAI22_X1 port map( A1 => n4660, A2 => n19307, B1 => n3779, B2 => 
                           n19301, ZN => n5506);
   U4373 : OAI22_X1 port map( A1 => n4659, A2 => n19108, B1 => n3778, B2 => 
                           n19102, ZN => n5457);
   U4374 : OAI22_X1 port map( A1 => n4659, A2 => n19307, B1 => n3778, B2 => 
                           n19301, ZN => n5437);
   U4375 : OAI22_X1 port map( A1 => n4658, A2 => n19108, B1 => n3777, B2 => 
                           n19102, ZN => n5389);
   U4376 : OAI22_X1 port map( A1 => n4658, A2 => n19307, B1 => n3777, B2 => 
                           n19301, ZN => n5369);
   U4377 : OAI22_X1 port map( A1 => n4580, A2 => n19080, B1 => n4511, B2 => 
                           n19074, ZN => n11659);
   U4378 : OAI22_X1 port map( A1 => n4580, A2 => n19279, B1 => n4511, B2 => 
                           n19273, ZN => n11620);
   U4379 : OAI22_X1 port map( A1 => n4579, A2 => n19080, B1 => n4510, B2 => 
                           n19074, ZN => n11533);
   U4380 : OAI22_X1 port map( A1 => n4579, A2 => n19279, B1 => n4510, B2 => 
                           n19273, ZN => n11515);
   U4381 : OAI22_X1 port map( A1 => n4578, A2 => n19080, B1 => n4509, B2 => 
                           n19074, ZN => n11466);
   U4382 : OAI22_X1 port map( A1 => n4578, A2 => n19279, B1 => n4509, B2 => 
                           n19273, ZN => n11448);
   U4383 : OAI22_X1 port map( A1 => n4577, A2 => n19080, B1 => n4508, B2 => 
                           n19074, ZN => n11399);
   U4384 : OAI22_X1 port map( A1 => n4577, A2 => n19279, B1 => n4508, B2 => 
                           n19273, ZN => n11380);
   U4385 : OAI22_X1 port map( A1 => n4576, A2 => n19080, B1 => n4507, B2 => 
                           n19074, ZN => n11332);
   U4386 : OAI22_X1 port map( A1 => n4576, A2 => n19279, B1 => n4507, B2 => 
                           n19273, ZN => n11313);
   U4387 : OAI22_X1 port map( A1 => n4575, A2 => n19080, B1 => n4506, B2 => 
                           n19074, ZN => n11264);
   U4388 : OAI22_X1 port map( A1 => n4575, A2 => n19279, B1 => n4506, B2 => 
                           n19273, ZN => n11246);
   U4389 : OAI22_X1 port map( A1 => n4574, A2 => n19080, B1 => n4505, B2 => 
                           n19074, ZN => n11197);
   U4390 : OAI22_X1 port map( A1 => n4574, A2 => n19279, B1 => n4505, B2 => 
                           n19273, ZN => n11179);
   U4391 : OAI22_X1 port map( A1 => n4573, A2 => n19080, B1 => n4504, B2 => 
                           n19074, ZN => n11130);
   U4392 : OAI22_X1 port map( A1 => n4573, A2 => n19279, B1 => n4504, B2 => 
                           n19273, ZN => n11111);
   U4393 : OAI22_X1 port map( A1 => n4572, A2 => n19080, B1 => n4503, B2 => 
                           n19074, ZN => n11062);
   U4394 : OAI22_X1 port map( A1 => n4572, A2 => n19279, B1 => n4503, B2 => 
                           n19273, ZN => n11044);
   U4395 : OAI22_X1 port map( A1 => n4571, A2 => n19080, B1 => n4502, B2 => 
                           n19074, ZN => n10995);
   U4396 : OAI22_X1 port map( A1 => n4571, A2 => n19279, B1 => n4502, B2 => 
                           n19273, ZN => n10977);
   U4397 : OAI22_X1 port map( A1 => n4570, A2 => n19080, B1 => n4501, B2 => 
                           n19074, ZN => n10928);
   U4398 : OAI22_X1 port map( A1 => n4570, A2 => n19279, B1 => n4501, B2 => 
                           n19273, ZN => n10910);
   U4399 : OAI22_X1 port map( A1 => n4569, A2 => n19080, B1 => n4500, B2 => 
                           n19074, ZN => n10861);
   U4400 : OAI22_X1 port map( A1 => n4569, A2 => n19279, B1 => n4500, B2 => 
                           n19273, ZN => n10842);
   U4401 : OAI22_X1 port map( A1 => n4568, A2 => n19081, B1 => n4499, B2 => 
                           n19075, ZN => n10793);
   U4402 : OAI22_X1 port map( A1 => n4568, A2 => n19280, B1 => n4499, B2 => 
                           n19274, ZN => n10775);
   U4403 : OAI22_X1 port map( A1 => n4567, A2 => n19081, B1 => n4498, B2 => 
                           n19075, ZN => n10726);
   U4404 : OAI22_X1 port map( A1 => n4567, A2 => n19280, B1 => n4498, B2 => 
                           n19274, ZN => n10708);
   U4405 : OAI22_X1 port map( A1 => n4566, A2 => n19081, B1 => n4497, B2 => 
                           n19075, ZN => n10659);
   U4406 : OAI22_X1 port map( A1 => n4566, A2 => n19280, B1 => n4497, B2 => 
                           n19274, ZN => n10640);
   U4407 : OAI22_X1 port map( A1 => n4565, A2 => n19081, B1 => n4496, B2 => 
                           n19075, ZN => n10592);
   U4408 : OAI22_X1 port map( A1 => n4565, A2 => n19280, B1 => n4496, B2 => 
                           n19274, ZN => n10573);
   U4409 : OAI22_X1 port map( A1 => n4564, A2 => n19081, B1 => n4495, B2 => 
                           n19075, ZN => n10524);
   U4410 : OAI22_X1 port map( A1 => n4564, A2 => n19280, B1 => n4495, B2 => 
                           n19274, ZN => n10506);
   U4411 : OAI22_X1 port map( A1 => n4563, A2 => n19081, B1 => n4494, B2 => 
                           n19075, ZN => n10457);
   U4412 : OAI22_X1 port map( A1 => n4563, A2 => n19280, B1 => n4494, B2 => 
                           n19274, ZN => n10439);
   U4413 : OAI22_X1 port map( A1 => n4562, A2 => n19081, B1 => n4493, B2 => 
                           n19075, ZN => n10390);
   U4414 : OAI22_X1 port map( A1 => n4562, A2 => n19280, B1 => n4493, B2 => 
                           n19274, ZN => n10371);
   U4415 : OAI22_X1 port map( A1 => n4561, A2 => n19081, B1 => n4492, B2 => 
                           n19075, ZN => n10322);
   U4416 : OAI22_X1 port map( A1 => n4561, A2 => n19280, B1 => n4492, B2 => 
                           n19274, ZN => n10304);
   U4417 : OAI22_X1 port map( A1 => n4560, A2 => n19081, B1 => n4491, B2 => 
                           n19075, ZN => n10255);
   U4418 : OAI22_X1 port map( A1 => n4560, A2 => n19280, B1 => n4491, B2 => 
                           n19274, ZN => n10237);
   U4419 : OAI22_X1 port map( A1 => n4559, A2 => n19081, B1 => n4490, B2 => 
                           n19075, ZN => n10188);
   U4420 : OAI22_X1 port map( A1 => n4559, A2 => n19280, B1 => n4490, B2 => 
                           n19274, ZN => n10170);
   U4421 : OAI22_X1 port map( A1 => n4558, A2 => n19081, B1 => n4489, B2 => 
                           n19075, ZN => n10121);
   U4422 : OAI22_X1 port map( A1 => n4558, A2 => n19280, B1 => n4489, B2 => 
                           n19274, ZN => n10102);
   U4423 : OAI22_X1 port map( A1 => n4557, A2 => n19081, B1 => n4488, B2 => 
                           n19075, ZN => n10053);
   U4424 : OAI22_X1 port map( A1 => n4557, A2 => n19280, B1 => n4488, B2 => 
                           n19274, ZN => n10035);
   U4425 : OAI22_X1 port map( A1 => n4556, A2 => n19082, B1 => n4487, B2 => 
                           n19076, ZN => n9986);
   U4426 : OAI22_X1 port map( A1 => n4556, A2 => n19281, B1 => n4487, B2 => 
                           n19275, ZN => n9968);
   U4427 : OAI22_X1 port map( A1 => n4555, A2 => n19082, B1 => n4486, B2 => 
                           n19076, ZN => n9919);
   U4428 : OAI22_X1 port map( A1 => n4555, A2 => n19281, B1 => n4486, B2 => 
                           n19275, ZN => n9900);
   U4429 : OAI22_X1 port map( A1 => n4554, A2 => n19082, B1 => n4485, B2 => 
                           n19076, ZN => n9852);
   U4430 : OAI22_X1 port map( A1 => n4554, A2 => n19281, B1 => n4485, B2 => 
                           n19275, ZN => n9833);
   U4431 : OAI22_X1 port map( A1 => n4553, A2 => n19082, B1 => n4484, B2 => 
                           n19076, ZN => n9784);
   U4432 : OAI22_X1 port map( A1 => n4553, A2 => n19281, B1 => n4484, B2 => 
                           n19275, ZN => n9766);
   U4433 : OAI22_X1 port map( A1 => n4552, A2 => n19082, B1 => n4483, B2 => 
                           n19076, ZN => n9717);
   U4434 : OAI22_X1 port map( A1 => n4552, A2 => n19281, B1 => n4483, B2 => 
                           n19275, ZN => n9699);
   U4435 : OAI22_X1 port map( A1 => n4551, A2 => n19082, B1 => n4482, B2 => 
                           n19076, ZN => n9650);
   U4436 : OAI22_X1 port map( A1 => n4551, A2 => n19281, B1 => n4482, B2 => 
                           n19275, ZN => n9631);
   U4437 : OAI22_X1 port map( A1 => n4550, A2 => n19082, B1 => n4481, B2 => 
                           n19076, ZN => n9582);
   U4438 : OAI22_X1 port map( A1 => n4550, A2 => n19281, B1 => n4481, B2 => 
                           n19275, ZN => n9564);
   U4439 : OAI22_X1 port map( A1 => n4549, A2 => n19082, B1 => n4480, B2 => 
                           n19076, ZN => n9515);
   U4440 : OAI22_X1 port map( A1 => n4549, A2 => n19281, B1 => n4480, B2 => 
                           n19275, ZN => n9497);
   U4441 : OAI22_X1 port map( A1 => n4548, A2 => n19082, B1 => n4479, B2 => 
                           n19076, ZN => n9448);
   U4442 : OAI22_X1 port map( A1 => n4548, A2 => n19281, B1 => n4479, B2 => 
                           n19275, ZN => n9430);
   U4443 : OAI22_X1 port map( A1 => n4547, A2 => n19082, B1 => n4478, B2 => 
                           n19076, ZN => n9381);
   U4444 : OAI22_X1 port map( A1 => n4547, A2 => n19281, B1 => n4478, B2 => 
                           n19275, ZN => n9362);
   U4445 : OAI22_X1 port map( A1 => n4546, A2 => n19082, B1 => n4477, B2 => 
                           n19076, ZN => n9313);
   U4446 : OAI22_X1 port map( A1 => n4546, A2 => n19281, B1 => n4477, B2 => 
                           n19275, ZN => n9295);
   U4447 : OAI22_X1 port map( A1 => n4545, A2 => n19082, B1 => n4476, B2 => 
                           n19076, ZN => n7006);
   U4448 : OAI22_X1 port map( A1 => n4545, A2 => n19281, B1 => n4476, B2 => 
                           n19275, ZN => n6988);
   U4449 : OAI22_X1 port map( A1 => n4544, A2 => n19083, B1 => n4475, B2 => 
                           n19077, ZN => n6939);
   U4450 : OAI22_X1 port map( A1 => n4544, A2 => n19282, B1 => n4475, B2 => 
                           n19276, ZN => n6921);
   U4451 : OAI22_X1 port map( A1 => n4543, A2 => n19083, B1 => n4474, B2 => 
                           n19077, ZN => n6873);
   U4452 : OAI22_X1 port map( A1 => n4543, A2 => n19282, B1 => n4474, B2 => 
                           n19276, ZN => n6854);
   U4453 : OAI22_X1 port map( A1 => n4542, A2 => n19083, B1 => n4473, B2 => 
                           n19077, ZN => n6806);
   U4454 : OAI22_X1 port map( A1 => n4542, A2 => n19282, B1 => n4473, B2 => 
                           n19276, ZN => n6787);
   U4455 : OAI22_X1 port map( A1 => n4541, A2 => n19083, B1 => n4472, B2 => 
                           n19077, ZN => n6738);
   U4456 : OAI22_X1 port map( A1 => n4541, A2 => n19282, B1 => n4472, B2 => 
                           n19276, ZN => n6720);
   U4457 : OAI22_X1 port map( A1 => n4540, A2 => n19083, B1 => n4471, B2 => 
                           n19077, ZN => n6671);
   U4458 : OAI22_X1 port map( A1 => n4540, A2 => n19282, B1 => n4471, B2 => 
                           n19276, ZN => n6653);
   U4459 : OAI22_X1 port map( A1 => n4539, A2 => n19083, B1 => n4470, B2 => 
                           n19077, ZN => n6604);
   U4460 : OAI22_X1 port map( A1 => n4539, A2 => n19282, B1 => n4470, B2 => 
                           n19276, ZN => n6586);
   U4461 : OAI22_X1 port map( A1 => n4538, A2 => n19083, B1 => n4469, B2 => 
                           n19077, ZN => n6538);
   U4462 : OAI22_X1 port map( A1 => n4538, A2 => n19282, B1 => n4469, B2 => 
                           n19276, ZN => n6520);
   U4463 : OAI22_X1 port map( A1 => n4537, A2 => n19083, B1 => n4468, B2 => 
                           n19077, ZN => n6472);
   U4464 : OAI22_X1 port map( A1 => n4537, A2 => n19282, B1 => n4468, B2 => 
                           n19276, ZN => n6454);
   U4465 : OAI22_X1 port map( A1 => n4536, A2 => n19083, B1 => n4467, B2 => 
                           n19077, ZN => n6406);
   U4466 : OAI22_X1 port map( A1 => n4536, A2 => n19282, B1 => n4467, B2 => 
                           n19276, ZN => n6388);
   U4467 : OAI22_X1 port map( A1 => n4535, A2 => n19083, B1 => n4466, B2 => 
                           n19077, ZN => n6340);
   U4468 : OAI22_X1 port map( A1 => n4535, A2 => n19282, B1 => n4466, B2 => 
                           n19276, ZN => n6322);
   U4469 : OAI22_X1 port map( A1 => n4534, A2 => n19083, B1 => n4465, B2 => 
                           n19077, ZN => n6274);
   U4470 : OAI22_X1 port map( A1 => n4534, A2 => n19282, B1 => n4465, B2 => 
                           n19276, ZN => n6256);
   U4471 : OAI22_X1 port map( A1 => n4533, A2 => n19083, B1 => n4464, B2 => 
                           n19077, ZN => n6208);
   U4472 : OAI22_X1 port map( A1 => n4533, A2 => n19282, B1 => n4464, B2 => 
                           n19276, ZN => n6190);
   U4473 : OAI22_X1 port map( A1 => n4532, A2 => n19084, B1 => n4463, B2 => 
                           n19078, ZN => n6142);
   U4474 : OAI22_X1 port map( A1 => n4532, A2 => n19283, B1 => n4463, B2 => 
                           n19277, ZN => n6124);
   U4475 : OAI22_X1 port map( A1 => n4531, A2 => n19084, B1 => n4462, B2 => 
                           n19078, ZN => n6076);
   U4476 : OAI22_X1 port map( A1 => n4531, A2 => n19283, B1 => n4462, B2 => 
                           n19277, ZN => n6058);
   U4477 : OAI22_X1 port map( A1 => n4530, A2 => n19084, B1 => n4461, B2 => 
                           n19078, ZN => n6008);
   U4478 : OAI22_X1 port map( A1 => n4530, A2 => n19283, B1 => n4461, B2 => 
                           n19277, ZN => n5990);
   U4479 : OAI22_X1 port map( A1 => n4529, A2 => n19084, B1 => n4460, B2 => 
                           n19078, ZN => n5940);
   U4480 : OAI22_X1 port map( A1 => n4529, A2 => n19283, B1 => n4460, B2 => 
                           n19277, ZN => n5922);
   U4481 : OAI22_X1 port map( A1 => n4528, A2 => n19084, B1 => n4459, B2 => 
                           n19078, ZN => n5873);
   U4482 : OAI22_X1 port map( A1 => n4528, A2 => n19283, B1 => n4459, B2 => 
                           n19277, ZN => n5855);
   U4483 : OAI22_X1 port map( A1 => n4527, A2 => n19084, B1 => n4458, B2 => 
                           n19078, ZN => n5806);
   U4484 : OAI22_X1 port map( A1 => n4527, A2 => n19283, B1 => n4458, B2 => 
                           n19277, ZN => n5788);
   U4485 : OAI22_X1 port map( A1 => n4526, A2 => n19084, B1 => n4457, B2 => 
                           n19078, ZN => n5734);
   U4486 : OAI22_X1 port map( A1 => n4526, A2 => n19283, B1 => n4457, B2 => 
                           n19277, ZN => n5716);
   U4487 : OAI22_X1 port map( A1 => n4525, A2 => n19084, B1 => n4456, B2 => 
                           n19078, ZN => n5664);
   U4488 : OAI22_X1 port map( A1 => n4525, A2 => n19283, B1 => n4456, B2 => 
                           n19277, ZN => n5646);
   U4489 : OAI22_X1 port map( A1 => n4524, A2 => n19084, B1 => n4455, B2 => 
                           n19078, ZN => n5596);
   U4490 : OAI22_X1 port map( A1 => n4524, A2 => n19283, B1 => n4455, B2 => 
                           n19277, ZN => n5578);
   U4491 : OAI22_X1 port map( A1 => n4523, A2 => n19084, B1 => n4454, B2 => 
                           n19078, ZN => n5527);
   U4492 : OAI22_X1 port map( A1 => n4523, A2 => n19283, B1 => n4454, B2 => 
                           n19277, ZN => n5509);
   U4493 : OAI22_X1 port map( A1 => n4522, A2 => n19084, B1 => n4453, B2 => 
                           n19078, ZN => n5458);
   U4494 : OAI22_X1 port map( A1 => n4522, A2 => n19283, B1 => n4453, B2 => 
                           n19277, ZN => n5440);
   U4495 : OAI22_X1 port map( A1 => n4521, A2 => n19084, B1 => n4452, B2 => 
                           n19078, ZN => n5390);
   U4496 : OAI22_X1 port map( A1 => n4521, A2 => n19283, B1 => n4452, B2 => 
                           n19277, ZN => n5372);
   U4497 : OAI22_X1 port map( A1 => n3577, A2 => n19151, B1 => n1733, B2 => 
                           n19145, ZN => n5316);
   U4498 : OAI22_X1 port map( A1 => n3577, A2 => n19350, B1 => n1733, B2 => 
                           n19344, ZN => n5296);
   U4499 : OAI22_X1 port map( A1 => n3576, A2 => n19151, B1 => n1732, B2 => 
                           n19145, ZN => n4447);
   U4500 : OAI22_X1 port map( A1 => n3576, A2 => n19350, B1 => n1732, B2 => 
                           n19344, ZN => n4107);
   U4501 : OAI22_X1 port map( A1 => n3575, A2 => n19151, B1 => n1731, B2 => 
                           n19145, ZN => n3290);
   U4502 : OAI22_X1 port map( A1 => n3575, A2 => n19350, B1 => n1731, B2 => 
                           n19344, ZN => n3250);
   U4503 : OAI22_X1 port map( A1 => n3574, A2 => n19151, B1 => n1730, B2 => 
                           n19145, ZN => n3117);
   U4504 : OAI22_X1 port map( A1 => n3574, A2 => n19350, B1 => n1730, B2 => 
                           n19344, ZN => n3000);
   U4505 : NAND2_X1 port map( A1 => cwp(1), A2 => n11753, ZN => n11739);
   U4506 : OAI22_X1 port map( A1 => n4542, A2 => n18927, B1 => n4745, B2 => 
                           n18921, ZN => n6825);
   U4507 : OAI22_X1 port map( A1 => n4541, A2 => n18927, B1 => n4744, B2 => 
                           n18921, ZN => n6758);
   U4508 : OAI22_X1 port map( A1 => n4540, A2 => n18927, B1 => n4743, B2 => 
                           n18921, ZN => n6690);
   U4509 : OAI22_X1 port map( A1 => n4539, A2 => n18927, B1 => n4742, B2 => 
                           n18921, ZN => n6623);
   U4510 : OAI22_X1 port map( A1 => n4538, A2 => n18927, B1 => n4741, B2 => 
                           n18921, ZN => n6557);
   U4511 : OAI22_X1 port map( A1 => n4537, A2 => n18927, B1 => n4740, B2 => 
                           n18921, ZN => n6491);
   U4512 : OAI22_X1 port map( A1 => n4536, A2 => n18927, B1 => n4739, B2 => 
                           n18921, ZN => n6425);
   U4513 : OAI22_X1 port map( A1 => n4535, A2 => n18927, B1 => n4738, B2 => 
                           n18921, ZN => n6359);
   U4514 : OAI22_X1 port map( A1 => n4534, A2 => n18927, B1 => n4737, B2 => 
                           n18921, ZN => n6293);
   U4515 : OAI22_X1 port map( A1 => n4533, A2 => n18927, B1 => n4736, B2 => 
                           n18921, ZN => n6227);
   U4516 : OAI22_X1 port map( A1 => n4532, A2 => n18928, B1 => n4735, B2 => 
                           n18922, ZN => n6161);
   U4517 : OAI22_X1 port map( A1 => n4531, A2 => n18928, B1 => n4734, B2 => 
                           n18922, ZN => n6095);
   U4518 : OAI22_X1 port map( A1 => n4530, A2 => n18928, B1 => n4733, B2 => 
                           n18922, ZN => n6027);
   U4519 : OAI22_X1 port map( A1 => n4529, A2 => n18928, B1 => n4732, B2 => 
                           n18922, ZN => n5959);
   U4520 : OAI22_X1 port map( A1 => n4528, A2 => n18928, B1 => n4731, B2 => 
                           n18922, ZN => n5892);
   U4521 : OAI22_X1 port map( A1 => n4527, A2 => n18928, B1 => n4730, B2 => 
                           n18922, ZN => n5825);
   U4522 : OAI22_X1 port map( A1 => n4526, A2 => n18928, B1 => n4729, B2 => 
                           n18922, ZN => n5753);
   U4523 : OAI22_X1 port map( A1 => n4525, A2 => n18928, B1 => n4728, B2 => 
                           n18922, ZN => n5683);
   U4524 : OAI22_X1 port map( A1 => n4524, A2 => n18928, B1 => n4727, B2 => 
                           n18922, ZN => n5615);
   U4525 : OAI22_X1 port map( A1 => n4523, A2 => n18928, B1 => n4726, B2 => 
                           n18922, ZN => n5546);
   U4526 : OAI22_X1 port map( A1 => n4522, A2 => n18928, B1 => n4725, B2 => 
                           n18922, ZN => n5477);
   U4527 : OAI22_X1 port map( A1 => n4521, A2 => n18928, B1 => n4724, B2 => 
                           n18922, ZN => n5409);
   U4528 : OAI22_X1 port map( A1 => n4580, A2 => n18924, B1 => n4783, B2 => 
                           n18918, ZN => n11714);
   U4529 : OAI22_X1 port map( A1 => n4579, A2 => n18924, B1 => n4782, B2 => 
                           n18918, ZN => n11553);
   U4530 : OAI22_X1 port map( A1 => n4578, A2 => n18924, B1 => n4781, B2 => 
                           n18918, ZN => n11485);
   U4531 : OAI22_X1 port map( A1 => n4577, A2 => n18924, B1 => n4780, B2 => 
                           n18918, ZN => n11418);
   U4532 : OAI22_X1 port map( A1 => n4576, A2 => n18924, B1 => n4779, B2 => 
                           n18918, ZN => n11351);
   U4533 : OAI22_X1 port map( A1 => n4575, A2 => n18924, B1 => n4778, B2 => 
                           n18918, ZN => n11284);
   U4534 : OAI22_X1 port map( A1 => n4574, A2 => n18924, B1 => n4777, B2 => 
                           n18918, ZN => n11216);
   U4535 : OAI22_X1 port map( A1 => n4573, A2 => n18924, B1 => n4776, B2 => 
                           n18918, ZN => n11149);
   U4536 : OAI22_X1 port map( A1 => n4572, A2 => n18924, B1 => n4775, B2 => 
                           n18918, ZN => n11082);
   U4537 : OAI22_X1 port map( A1 => n4571, A2 => n18924, B1 => n4774, B2 => 
                           n18918, ZN => n11015);
   U4538 : OAI22_X1 port map( A1 => n4570, A2 => n18924, B1 => n4773, B2 => 
                           n18918, ZN => n10947);
   U4539 : OAI22_X1 port map( A1 => n4569, A2 => n18924, B1 => n4772, B2 => 
                           n18918, ZN => n10880);
   U4540 : OAI22_X1 port map( A1 => n4568, A2 => n18925, B1 => n4771, B2 => 
                           n18919, ZN => n10813);
   U4541 : OAI22_X1 port map( A1 => n4567, A2 => n18925, B1 => n4770, B2 => 
                           n18919, ZN => n10745);
   U4542 : OAI22_X1 port map( A1 => n4566, A2 => n18925, B1 => n4769, B2 => 
                           n18919, ZN => n10678);
   U4543 : OAI22_X1 port map( A1 => n4565, A2 => n18925, B1 => n4768, B2 => 
                           n18919, ZN => n10611);
   U4544 : OAI22_X1 port map( A1 => n4564, A2 => n18925, B1 => n4767, B2 => 
                           n18919, ZN => n10544);
   U4545 : OAI22_X1 port map( A1 => n4563, A2 => n18925, B1 => n4766, B2 => 
                           n18919, ZN => n10476);
   U4546 : OAI22_X1 port map( A1 => n4562, A2 => n18925, B1 => n4765, B2 => 
                           n18919, ZN => n10409);
   U4547 : OAI22_X1 port map( A1 => n4561, A2 => n18925, B1 => n4764, B2 => 
                           n18919, ZN => n10342);
   U4548 : OAI22_X1 port map( A1 => n4560, A2 => n18925, B1 => n4763, B2 => 
                           n18919, ZN => n10275);
   U4549 : OAI22_X1 port map( A1 => n4559, A2 => n18925, B1 => n4762, B2 => 
                           n18919, ZN => n10207);
   U4550 : OAI22_X1 port map( A1 => n4558, A2 => n18925, B1 => n4761, B2 => 
                           n18919, ZN => n10140);
   U4551 : OAI22_X1 port map( A1 => n4557, A2 => n18925, B1 => n4760, B2 => 
                           n18919, ZN => n10073);
   U4552 : OAI22_X1 port map( A1 => n4556, A2 => n18926, B1 => n4759, B2 => 
                           n18920, ZN => n10005);
   U4553 : OAI22_X1 port map( A1 => n4555, A2 => n18926, B1 => n4758, B2 => 
                           n18920, ZN => n9938);
   U4554 : OAI22_X1 port map( A1 => n4554, A2 => n18926, B1 => n4757, B2 => 
                           n18920, ZN => n9871);
   U4555 : OAI22_X1 port map( A1 => n4553, A2 => n18926, B1 => n4756, B2 => 
                           n18920, ZN => n9804);
   U4556 : OAI22_X1 port map( A1 => n4552, A2 => n18926, B1 => n4755, B2 => 
                           n18920, ZN => n9736);
   U4557 : OAI22_X1 port map( A1 => n4551, A2 => n18926, B1 => n4754, B2 => 
                           n18920, ZN => n9669);
   U4558 : OAI22_X1 port map( A1 => n4550, A2 => n18926, B1 => n4753, B2 => 
                           n18920, ZN => n9602);
   U4559 : OAI22_X1 port map( A1 => n4549, A2 => n18926, B1 => n4752, B2 => 
                           n18920, ZN => n9535);
   U4560 : OAI22_X1 port map( A1 => n4548, A2 => n18926, B1 => n4751, B2 => 
                           n18920, ZN => n9467);
   U4561 : OAI22_X1 port map( A1 => n4547, A2 => n18926, B1 => n4750, B2 => 
                           n18920, ZN => n9400);
   U4562 : OAI22_X1 port map( A1 => n4546, A2 => n18926, B1 => n4749, B2 => 
                           n18920, ZN => n9333);
   U4563 : OAI22_X1 port map( A1 => n4545, A2 => n18926, B1 => n4748, B2 => 
                           n18920, ZN => n9266);
   U4564 : OAI22_X1 port map( A1 => n4544, A2 => n18927, B1 => n4747, B2 => 
                           n18921, ZN => n6959);
   U4565 : OAI22_X1 port map( A1 => n4543, A2 => n18927, B1 => n4746, B2 => 
                           n18921, ZN => n6892);
   U4566 : OAI22_X1 port map( A1 => n4948, A2 => n18975, B1 => n5014, B2 => 
                           n18969, ZN => n6753);
   U4567 : OAI22_X1 port map( A1 => n4947, A2 => n18975, B1 => n5013, B2 => 
                           n18969, ZN => n6685);
   U4568 : OAI22_X1 port map( A1 => n4946, A2 => n18975, B1 => n5012, B2 => 
                           n18969, ZN => n6618);
   U4569 : OAI22_X1 port map( A1 => n4945, A2 => n18975, B1 => n5011, B2 => 
                           n18969, ZN => n6552);
   U4570 : OAI22_X1 port map( A1 => n4944, A2 => n18975, B1 => n5010, B2 => 
                           n18969, ZN => n6486);
   U4571 : OAI22_X1 port map( A1 => n4943, A2 => n18975, B1 => n5009, B2 => 
                           n18969, ZN => n6420);
   U4572 : OAI22_X1 port map( A1 => n4942, A2 => n18975, B1 => n5008, B2 => 
                           n18969, ZN => n6354);
   U4573 : OAI22_X1 port map( A1 => n4941, A2 => n18975, B1 => n5007, B2 => 
                           n18969, ZN => n6288);
   U4574 : OAI22_X1 port map( A1 => n4940, A2 => n18975, B1 => n5006, B2 => 
                           n18969, ZN => n6222);
   U4575 : OAI22_X1 port map( A1 => n4975, A2 => n18973, B1 => n5041, B2 => 
                           n18967, ZN => n10808);
   U4576 : OAI22_X1 port map( A1 => n4974, A2 => n18973, B1 => n5040, B2 => 
                           n18967, ZN => n10740);
   U4577 : OAI22_X1 port map( A1 => n4973, A2 => n18973, B1 => n5039, B2 => 
                           n18967, ZN => n10673);
   U4578 : OAI22_X1 port map( A1 => n4972, A2 => n18973, B1 => n5038, B2 => 
                           n18967, ZN => n10606);
   U4579 : OAI22_X1 port map( A1 => n4971, A2 => n18973, B1 => n5037, B2 => 
                           n18967, ZN => n10539);
   U4580 : OAI22_X1 port map( A1 => n4970, A2 => n18973, B1 => n5036, B2 => 
                           n18967, ZN => n10471);
   U4581 : OAI22_X1 port map( A1 => n4969, A2 => n18973, B1 => n5035, B2 => 
                           n18967, ZN => n10404);
   U4582 : OAI22_X1 port map( A1 => n4968, A2 => n18973, B1 => n5034, B2 => 
                           n18967, ZN => n10337);
   U4583 : OAI22_X1 port map( A1 => n4967, A2 => n18973, B1 => n5033, B2 => 
                           n18967, ZN => n10269);
   U4584 : OAI22_X1 port map( A1 => n4966, A2 => n18973, B1 => n5032, B2 => 
                           n18967, ZN => n10202);
   U4585 : OAI22_X1 port map( A1 => n4965, A2 => n18973, B1 => n5031, B2 => 
                           n18967, ZN => n10135);
   U4586 : OAI22_X1 port map( A1 => n4964, A2 => n18973, B1 => n5030, B2 => 
                           n18967, ZN => n10068);
   U4587 : OAI22_X1 port map( A1 => n4963, A2 => n18974, B1 => n5029, B2 => 
                           n18968, ZN => n10000);
   U4588 : OAI22_X1 port map( A1 => n4962, A2 => n18974, B1 => n5028, B2 => 
                           n18968, ZN => n9933);
   U4589 : OAI22_X1 port map( A1 => n4961, A2 => n18974, B1 => n5027, B2 => 
                           n18968, ZN => n9866);
   U4590 : OAI22_X1 port map( A1 => n4960, A2 => n18974, B1 => n5026, B2 => 
                           n18968, ZN => n9799);
   U4591 : OAI22_X1 port map( A1 => n4959, A2 => n18974, B1 => n5025, B2 => 
                           n18968, ZN => n9731);
   U4592 : OAI22_X1 port map( A1 => n4958, A2 => n18974, B1 => n5024, B2 => 
                           n18968, ZN => n9664);
   U4593 : OAI22_X1 port map( A1 => n4957, A2 => n18974, B1 => n5023, B2 => 
                           n18968, ZN => n9597);
   U4594 : OAI22_X1 port map( A1 => n4956, A2 => n18974, B1 => n5022, B2 => 
                           n18968, ZN => n9529);
   U4595 : OAI22_X1 port map( A1 => n4955, A2 => n18974, B1 => n5021, B2 => 
                           n18968, ZN => n9462);
   U4596 : OAI22_X1 port map( A1 => n4954, A2 => n18974, B1 => n5020, B2 => 
                           n18968, ZN => n9395);
   U4597 : OAI22_X1 port map( A1 => n4953, A2 => n18974, B1 => n5019, B2 => 
                           n18968, ZN => n9328);
   U4598 : OAI22_X1 port map( A1 => n4952, A2 => n18974, B1 => n5018, B2 => 
                           n18968, ZN => n7020);
   U4599 : OAI22_X1 port map( A1 => n4951, A2 => n18975, B1 => n5017, B2 => 
                           n18969, ZN => n6954);
   U4600 : OAI22_X1 port map( A1 => n4950, A2 => n18975, B1 => n5016, B2 => 
                           n18969, ZN => n6887);
   U4601 : OAI22_X1 port map( A1 => n4939, A2 => n18976, B1 => n5005, B2 => 
                           n18970, ZN => n6156);
   U4602 : OAI22_X1 port map( A1 => n4938, A2 => n18976, B1 => n5004, B2 => 
                           n18970, ZN => n6090);
   U4603 : OAI22_X1 port map( A1 => n4937, A2 => n18976, B1 => n5003, B2 => 
                           n18970, ZN => n6022);
   U4604 : OAI22_X1 port map( A1 => n4936, A2 => n18976, B1 => n5002, B2 => 
                           n18970, ZN => n5954);
   U4605 : OAI22_X1 port map( A1 => n4935, A2 => n18976, B1 => n5001, B2 => 
                           n18970, ZN => n5887);
   U4606 : OAI22_X1 port map( A1 => n4934, A2 => n18976, B1 => n5000, B2 => 
                           n18970, ZN => n5820);
   U4607 : OAI22_X1 port map( A1 => n4933, A2 => n18976, B1 => n4999, B2 => 
                           n18970, ZN => n5748);
   U4608 : OAI22_X1 port map( A1 => n4932, A2 => n18976, B1 => n4998, B2 => 
                           n18970, ZN => n5678);
   U4609 : OAI22_X1 port map( A1 => n4931, A2 => n18976, B1 => n4997, B2 => 
                           n18970, ZN => n5610);
   U4610 : OAI22_X1 port map( A1 => n4930, A2 => n18976, B1 => n4996, B2 => 
                           n18970, ZN => n5541);
   U4611 : OAI22_X1 port map( A1 => n4929, A2 => n18976, B1 => n4995, B2 => 
                           n18970, ZN => n5472);
   U4612 : OAI22_X1 port map( A1 => n4928, A2 => n18976, B1 => n4994, B2 => 
                           n18970, ZN => n5404);
   U4613 : OAI22_X1 port map( A1 => n3637, A2 => n19146, B1 => n1796, B2 => 
                           n19140, ZN => n11649);
   U4614 : OAI22_X1 port map( A1 => n3637, A2 => n19345, B1 => n1796, B2 => 
                           n19339, ZN => n11608);
   U4615 : OAI22_X1 port map( A1 => n3636, A2 => n19146, B1 => n1795, B2 => 
                           n19140, ZN => n11529);
   U4616 : OAI22_X1 port map( A1 => n3636, A2 => n19345, B1 => n1795, B2 => 
                           n19339, ZN => n11509);
   U4617 : OAI22_X1 port map( A1 => n3635, A2 => n19146, B1 => n1794, B2 => 
                           n19140, ZN => n11462);
   U4618 : OAI22_X1 port map( A1 => n3635, A2 => n19345, B1 => n1794, B2 => 
                           n19339, ZN => n11442);
   U4619 : OAI22_X1 port map( A1 => n3634, A2 => n19146, B1 => n1793, B2 => 
                           n19140, ZN => n11395);
   U4620 : OAI22_X1 port map( A1 => n3634, A2 => n19345, B1 => n1793, B2 => 
                           n19339, ZN => n11374);
   U4621 : OAI22_X1 port map( A1 => n3633, A2 => n19146, B1 => n1792, B2 => 
                           n19140, ZN => n11327);
   U4622 : OAI22_X1 port map( A1 => n3633, A2 => n19345, B1 => n1792, B2 => 
                           n19339, ZN => n11307);
   U4623 : OAI22_X1 port map( A1 => n3632, A2 => n19146, B1 => n1791, B2 => 
                           n19140, ZN => n11260);
   U4624 : OAI22_X1 port map( A1 => n3632, A2 => n19345, B1 => n1791, B2 => 
                           n19339, ZN => n11240);
   U4625 : OAI22_X1 port map( A1 => n3631, A2 => n19146, B1 => n1790, B2 => 
                           n19140, ZN => n11193);
   U4626 : OAI22_X1 port map( A1 => n3631, A2 => n19345, B1 => n1790, B2 => 
                           n19339, ZN => n11173);
   U4627 : OAI22_X1 port map( A1 => n3630, A2 => n19146, B1 => n1789, B2 => 
                           n19140, ZN => n11126);
   U4628 : OAI22_X1 port map( A1 => n3630, A2 => n19345, B1 => n1789, B2 => 
                           n19339, ZN => n11105);
   U4629 : OAI22_X1 port map( A1 => n3629, A2 => n19146, B1 => n1788, B2 => 
                           n19140, ZN => n11058);
   U4630 : OAI22_X1 port map( A1 => n3629, A2 => n19345, B1 => n1788, B2 => 
                           n19339, ZN => n11038);
   U4631 : OAI22_X1 port map( A1 => n3628, A2 => n19146, B1 => n1787, B2 => 
                           n19140, ZN => n10991);
   U4632 : OAI22_X1 port map( A1 => n3628, A2 => n19345, B1 => n1787, B2 => 
                           n19339, ZN => n10971);
   U4633 : OAI22_X1 port map( A1 => n3627, A2 => n19146, B1 => n1786, B2 => 
                           n19140, ZN => n10924);
   U4634 : OAI22_X1 port map( A1 => n3627, A2 => n19345, B1 => n1786, B2 => 
                           n19339, ZN => n10903);
   U4635 : OAI22_X1 port map( A1 => n3626, A2 => n19146, B1 => n1785, B2 => 
                           n19140, ZN => n10857);
   U4636 : OAI22_X1 port map( A1 => n3626, A2 => n19345, B1 => n1785, B2 => 
                           n19339, ZN => n10836);
   U4637 : OAI22_X1 port map( A1 => n3625, A2 => n19147, B1 => n1784, B2 => 
                           n19141, ZN => n10789);
   U4638 : OAI22_X1 port map( A1 => n3625, A2 => n19346, B1 => n1784, B2 => 
                           n19340, ZN => n10769);
   U4639 : OAI22_X1 port map( A1 => n3624, A2 => n19147, B1 => n1783, B2 => 
                           n19141, ZN => n10722);
   U4640 : OAI22_X1 port map( A1 => n3624, A2 => n19346, B1 => n1783, B2 => 
                           n19340, ZN => n10702);
   U4641 : OAI22_X1 port map( A1 => n3623, A2 => n19147, B1 => n1782, B2 => 
                           n19141, ZN => n10655);
   U4642 : OAI22_X1 port map( A1 => n3623, A2 => n19346, B1 => n1782, B2 => 
                           n19340, ZN => n10634);
   U4643 : OAI22_X1 port map( A1 => n3622, A2 => n19147, B1 => n1781, B2 => 
                           n19141, ZN => n10587);
   U4644 : OAI22_X1 port map( A1 => n3622, A2 => n19346, B1 => n1781, B2 => 
                           n19340, ZN => n10567);
   U4645 : OAI22_X1 port map( A1 => n3621, A2 => n19147, B1 => n1780, B2 => 
                           n19141, ZN => n10520);
   U4646 : OAI22_X1 port map( A1 => n3621, A2 => n19346, B1 => n1780, B2 => 
                           n19340, ZN => n10500);
   U4647 : OAI22_X1 port map( A1 => n3620, A2 => n19147, B1 => n1779, B2 => 
                           n19141, ZN => n10453);
   U4648 : OAI22_X1 port map( A1 => n3620, A2 => n19346, B1 => n1779, B2 => 
                           n19340, ZN => n10433);
   U4649 : OAI22_X1 port map( A1 => n3619, A2 => n19147, B1 => n1778, B2 => 
                           n19141, ZN => n10386);
   U4650 : OAI22_X1 port map( A1 => n3619, A2 => n19346, B1 => n1778, B2 => 
                           n19340, ZN => n10365);
   U4651 : OAI22_X1 port map( A1 => n3618, A2 => n19147, B1 => n1777, B2 => 
                           n19141, ZN => n10318);
   U4652 : OAI22_X1 port map( A1 => n3618, A2 => n19346, B1 => n1777, B2 => 
                           n19340, ZN => n10298);
   U4653 : OAI22_X1 port map( A1 => n3617, A2 => n19147, B1 => n1776, B2 => 
                           n19141, ZN => n10251);
   U4654 : OAI22_X1 port map( A1 => n3617, A2 => n19346, B1 => n1776, B2 => 
                           n19340, ZN => n10231);
   U4655 : OAI22_X1 port map( A1 => n3616, A2 => n19147, B1 => n1775, B2 => 
                           n19141, ZN => n10184);
   U4656 : OAI22_X1 port map( A1 => n3616, A2 => n19346, B1 => n1775, B2 => 
                           n19340, ZN => n10163);
   U4657 : OAI22_X1 port map( A1 => n3615, A2 => n19147, B1 => n1774, B2 => 
                           n19141, ZN => n10117);
   U4658 : OAI22_X1 port map( A1 => n3615, A2 => n19346, B1 => n1774, B2 => 
                           n19340, ZN => n10096);
   U4659 : OAI22_X1 port map( A1 => n3614, A2 => n19147, B1 => n1773, B2 => 
                           n19141, ZN => n10049);
   U4660 : OAI22_X1 port map( A1 => n3614, A2 => n19346, B1 => n1773, B2 => 
                           n19340, ZN => n10029);
   U4661 : OAI22_X1 port map( A1 => n3613, A2 => n19148, B1 => n1772, B2 => 
                           n19142, ZN => n9982);
   U4662 : OAI22_X1 port map( A1 => n3613, A2 => n19347, B1 => n1772, B2 => 
                           n19341, ZN => n9962);
   U4663 : OAI22_X1 port map( A1 => n3612, A2 => n19148, B1 => n1771, B2 => 
                           n19142, ZN => n9915);
   U4664 : OAI22_X1 port map( A1 => n3612, A2 => n19347, B1 => n1771, B2 => 
                           n19341, ZN => n9894);
   U4665 : OAI22_X1 port map( A1 => n3611, A2 => n19148, B1 => n1770, B2 => 
                           n19142, ZN => n9847);
   U4666 : OAI22_X1 port map( A1 => n3611, A2 => n19347, B1 => n1770, B2 => 
                           n19341, ZN => n9827);
   U4667 : OAI22_X1 port map( A1 => n3610, A2 => n19148, B1 => n1769, B2 => 
                           n19142, ZN => n9780);
   U4668 : OAI22_X1 port map( A1 => n3610, A2 => n19347, B1 => n1769, B2 => 
                           n19341, ZN => n9760);
   U4669 : OAI22_X1 port map( A1 => n3609, A2 => n19148, B1 => n1768, B2 => 
                           n19142, ZN => n9713);
   U4670 : OAI22_X1 port map( A1 => n3609, A2 => n19347, B1 => n1768, B2 => 
                           n19341, ZN => n9693);
   U4671 : OAI22_X1 port map( A1 => n3608, A2 => n19148, B1 => n1767, B2 => 
                           n19142, ZN => n9646);
   U4672 : OAI22_X1 port map( A1 => n3608, A2 => n19347, B1 => n1767, B2 => 
                           n19341, ZN => n9625);
   U4673 : OAI22_X1 port map( A1 => n3607, A2 => n19148, B1 => n1766, B2 => 
                           n19142, ZN => n9578);
   U4674 : OAI22_X1 port map( A1 => n3607, A2 => n19347, B1 => n1766, B2 => 
                           n19341, ZN => n9558);
   U4675 : OAI22_X1 port map( A1 => n3606, A2 => n19148, B1 => n1765, B2 => 
                           n19142, ZN => n9511);
   U4676 : OAI22_X1 port map( A1 => n3606, A2 => n19347, B1 => n1765, B2 => 
                           n19341, ZN => n9491);
   U4677 : OAI22_X1 port map( A1 => n3605, A2 => n19148, B1 => n1764, B2 => 
                           n19142, ZN => n9444);
   U4678 : OAI22_X1 port map( A1 => n3605, A2 => n19347, B1 => n1764, B2 => 
                           n19341, ZN => n9423);
   U4679 : OAI22_X1 port map( A1 => n3604, A2 => n19148, B1 => n1763, B2 => 
                           n19142, ZN => n9377);
   U4680 : OAI22_X1 port map( A1 => n3604, A2 => n19347, B1 => n1763, B2 => 
                           n19341, ZN => n9356);
   U4681 : OAI22_X1 port map( A1 => n3603, A2 => n19148, B1 => n1762, B2 => 
                           n19142, ZN => n9309);
   U4682 : OAI22_X1 port map( A1 => n3603, A2 => n19347, B1 => n1762, B2 => 
                           n19341, ZN => n9289);
   U4683 : OAI22_X1 port map( A1 => n3602, A2 => n19148, B1 => n1761, B2 => 
                           n19142, ZN => n7002);
   U4684 : OAI22_X1 port map( A1 => n3602, A2 => n19347, B1 => n1761, B2 => 
                           n19341, ZN => n6982);
   U4685 : OAI22_X1 port map( A1 => n3601, A2 => n19149, B1 => n1760, B2 => 
                           n19143, ZN => n6935);
   U4686 : OAI22_X1 port map( A1 => n3601, A2 => n19348, B1 => n1760, B2 => 
                           n19342, ZN => n6915);
   U4687 : OAI22_X1 port map( A1 => n3600, A2 => n19149, B1 => n1759, B2 => 
                           n19143, ZN => n6869);
   U4688 : OAI22_X1 port map( A1 => n3600, A2 => n19348, B1 => n1759, B2 => 
                           n19342, ZN => n6848);
   U4689 : OAI22_X1 port map( A1 => n3599, A2 => n19149, B1 => n1758, B2 => 
                           n19143, ZN => n6801);
   U4690 : OAI22_X1 port map( A1 => n3599, A2 => n19348, B1 => n1758, B2 => 
                           n19342, ZN => n6781);
   U4691 : OAI22_X1 port map( A1 => n3598, A2 => n19149, B1 => n1757, B2 => 
                           n19143, ZN => n6734);
   U4692 : OAI22_X1 port map( A1 => n3598, A2 => n19348, B1 => n1757, B2 => 
                           n19342, ZN => n6714);
   U4693 : OAI22_X1 port map( A1 => n3597, A2 => n19149, B1 => n1756, B2 => 
                           n19143, ZN => n6667);
   U4694 : OAI22_X1 port map( A1 => n3597, A2 => n19348, B1 => n1756, B2 => 
                           n19342, ZN => n6647);
   U4695 : OAI22_X1 port map( A1 => n3596, A2 => n19149, B1 => n1755, B2 => 
                           n19143, ZN => n6600);
   U4696 : OAI22_X1 port map( A1 => n3596, A2 => n19348, B1 => n1755, B2 => 
                           n19342, ZN => n6580);
   U4697 : OAI22_X1 port map( A1 => n3595, A2 => n19149, B1 => n1754, B2 => 
                           n19143, ZN => n6534);
   U4698 : OAI22_X1 port map( A1 => n3595, A2 => n19348, B1 => n1754, B2 => 
                           n19342, ZN => n6514);
   U4699 : OAI22_X1 port map( A1 => n3594, A2 => n19149, B1 => n1753, B2 => 
                           n19143, ZN => n6468);
   U4700 : OAI22_X1 port map( A1 => n3594, A2 => n19348, B1 => n1753, B2 => 
                           n19342, ZN => n6448);
   U4701 : OAI22_X1 port map( A1 => n3593, A2 => n19149, B1 => n1752, B2 => 
                           n19143, ZN => n6402);
   U4702 : OAI22_X1 port map( A1 => n3593, A2 => n19348, B1 => n1752, B2 => 
                           n19342, ZN => n6382);
   U4703 : OAI22_X1 port map( A1 => n3592, A2 => n19149, B1 => n1751, B2 => 
                           n19143, ZN => n6336);
   U4704 : OAI22_X1 port map( A1 => n3592, A2 => n19348, B1 => n1751, B2 => 
                           n19342, ZN => n6316);
   U4705 : OAI22_X1 port map( A1 => n3591, A2 => n19149, B1 => n1750, B2 => 
                           n19143, ZN => n6270);
   U4706 : OAI22_X1 port map( A1 => n3591, A2 => n19348, B1 => n1750, B2 => 
                           n19342, ZN => n6250);
   U4707 : OAI22_X1 port map( A1 => n3590, A2 => n19149, B1 => n1749, B2 => 
                           n19143, ZN => n6204);
   U4708 : OAI22_X1 port map( A1 => n3590, A2 => n19348, B1 => n1749, B2 => 
                           n19342, ZN => n6184);
   U4709 : OAI22_X1 port map( A1 => n3589, A2 => n19150, B1 => n1745, B2 => 
                           n19144, ZN => n6138);
   U4710 : OAI22_X1 port map( A1 => n3589, A2 => n19349, B1 => n1745, B2 => 
                           n19343, ZN => n6118);
   U4711 : OAI22_X1 port map( A1 => n3588, A2 => n19150, B1 => n1744, B2 => 
                           n19144, ZN => n6072);
   U4712 : OAI22_X1 port map( A1 => n3588, A2 => n19349, B1 => n1744, B2 => 
                           n19343, ZN => n6052);
   U4713 : OAI22_X1 port map( A1 => n3587, A2 => n19150, B1 => n1743, B2 => 
                           n19144, ZN => n6004);
   U4714 : OAI22_X1 port map( A1 => n3587, A2 => n19349, B1 => n1743, B2 => 
                           n19343, ZN => n5984);
   U4715 : OAI22_X1 port map( A1 => n3586, A2 => n19150, B1 => n1742, B2 => 
                           n19144, ZN => n5936);
   U4716 : OAI22_X1 port map( A1 => n3586, A2 => n19349, B1 => n1742, B2 => 
                           n19343, ZN => n5916);
   U4717 : OAI22_X1 port map( A1 => n3585, A2 => n19150, B1 => n1741, B2 => 
                           n19144, ZN => n5869);
   U4718 : OAI22_X1 port map( A1 => n3585, A2 => n19349, B1 => n1741, B2 => 
                           n19343, ZN => n5849);
   U4719 : OAI22_X1 port map( A1 => n3584, A2 => n19150, B1 => n1740, B2 => 
                           n19144, ZN => n5802);
   U4720 : OAI22_X1 port map( A1 => n3584, A2 => n19349, B1 => n1740, B2 => 
                           n19343, ZN => n5782);
   U4721 : OAI22_X1 port map( A1 => n3583, A2 => n19150, B1 => n1739, B2 => 
                           n19144, ZN => n5730);
   U4722 : OAI22_X1 port map( A1 => n3583, A2 => n19349, B1 => n1739, B2 => 
                           n19343, ZN => n5710);
   U4723 : OAI22_X1 port map( A1 => n3582, A2 => n19150, B1 => n1738, B2 => 
                           n19144, ZN => n5660);
   U4724 : OAI22_X1 port map( A1 => n3582, A2 => n19349, B1 => n1738, B2 => 
                           n19343, ZN => n5640);
   U4725 : OAI22_X1 port map( A1 => n3581, A2 => n19150, B1 => n1737, B2 => 
                           n19144, ZN => n5592);
   U4726 : OAI22_X1 port map( A1 => n3581, A2 => n19349, B1 => n1737, B2 => 
                           n19343, ZN => n5572);
   U4727 : OAI22_X1 port map( A1 => n3580, A2 => n19150, B1 => n1736, B2 => 
                           n19144, ZN => n5523);
   U4728 : OAI22_X1 port map( A1 => n3580, A2 => n19349, B1 => n1736, B2 => 
                           n19343, ZN => n5503);
   U4729 : OAI22_X1 port map( A1 => n3579, A2 => n19150, B1 => n1735, B2 => 
                           n19144, ZN => n5454);
   U4730 : OAI22_X1 port map( A1 => n3579, A2 => n19349, B1 => n1735, B2 => 
                           n19343, ZN => n5434);
   U4731 : OAI22_X1 port map( A1 => n3578, A2 => n19150, B1 => n1734, B2 => 
                           n19144, ZN => n5386);
   U4732 : OAI22_X1 port map( A1 => n3578, A2 => n19349, B1 => n1734, B2 => 
                           n19343, ZN => n5366);
   U4733 : OAI22_X1 port map( A1 => n20367, A2 => n19690, B1 => n4917, B2 => 
                           n19705, ZN => n7667);
   U4734 : OAI22_X1 port map( A1 => n20370, A2 => n19690, B1 => n4916, B2 => 
                           n19705, ZN => n7668);
   U4735 : OAI22_X1 port map( A1 => n20373, A2 => n19690, B1 => n4915, B2 => 
                           n19705, ZN => n7669);
   U4736 : OAI22_X1 port map( A1 => n20376, A2 => n19690, B1 => n4914, B2 => 
                           n19705, ZN => n7670);
   U4737 : OAI22_X1 port map( A1 => n20379, A2 => n19690, B1 => n4913, B2 => 
                           n19704, ZN => n7671);
   U4738 : OAI22_X1 port map( A1 => n20382, A2 => n19690, B1 => n4912, B2 => 
                           n19704, ZN => n7672);
   U4739 : OAI22_X1 port map( A1 => n20385, A2 => n19690, B1 => n4911, B2 => 
                           n19704, ZN => n7673);
   U4740 : OAI22_X1 port map( A1 => n20388, A2 => n19690, B1 => n4910, B2 => 
                           n19704, ZN => n7674);
   U4741 : OAI22_X1 port map( A1 => n20391, A2 => n19690, B1 => n4909, B2 => 
                           n19703, ZN => n7675);
   U4742 : OAI22_X1 port map( A1 => n20394, A2 => n19690, B1 => n4908, B2 => 
                           n19703, ZN => n7676);
   U4743 : OAI22_X1 port map( A1 => n20397, A2 => n19690, B1 => n4907, B2 => 
                           n19703, ZN => n7677);
   U4744 : OAI22_X1 port map( A1 => n20400, A2 => n19690, B1 => n4906, B2 => 
                           n19703, ZN => n7678);
   U4745 : OAI22_X1 port map( A1 => n20403, A2 => n19689, B1 => n4905, B2 => 
                           n19702, ZN => n7679);
   U4746 : OAI22_X1 port map( A1 => n20406, A2 => n19689, B1 => n4904, B2 => 
                           n19702, ZN => n7680);
   U4747 : OAI22_X1 port map( A1 => n20409, A2 => n19689, B1 => n4903, B2 => 
                           n19702, ZN => n7681);
   U4748 : OAI22_X1 port map( A1 => n20412, A2 => n19689, B1 => n4902, B2 => 
                           n19702, ZN => n7682);
   U4749 : OAI22_X1 port map( A1 => n20415, A2 => n19689, B1 => n4901, B2 => 
                           n19701, ZN => n7683);
   U4750 : OAI22_X1 port map( A1 => n20418, A2 => n19689, B1 => n4900, B2 => 
                           n19701, ZN => n7684);
   U4751 : OAI22_X1 port map( A1 => n20421, A2 => n19689, B1 => n4899, B2 => 
                           n19701, ZN => n7685);
   U4752 : OAI22_X1 port map( A1 => n20424, A2 => n19689, B1 => n4898, B2 => 
                           n19701, ZN => n7686);
   U4753 : OAI22_X1 port map( A1 => n20427, A2 => n19689, B1 => n4897, B2 => 
                           n19700, ZN => n7687);
   U4754 : OAI22_X1 port map( A1 => n20430, A2 => n19689, B1 => n4896, B2 => 
                           n19700, ZN => n7688);
   U4755 : OAI22_X1 port map( A1 => n20433, A2 => n19689, B1 => n4895, B2 => 
                           n19700, ZN => n7689);
   U4756 : OAI22_X1 port map( A1 => n20436, A2 => n19689, B1 => n4894, B2 => 
                           n19700, ZN => n7690);
   U4757 : OAI22_X1 port map( A1 => n20439, A2 => n19688, B1 => n4893, B2 => 
                           n19699, ZN => n7691);
   U4758 : OAI22_X1 port map( A1 => n20442, A2 => n19688, B1 => n4892, B2 => 
                           n19699, ZN => n7692);
   U4759 : OAI22_X1 port map( A1 => n20445, A2 => n19688, B1 => n4891, B2 => 
                           n19699, ZN => n7693);
   U4760 : OAI22_X1 port map( A1 => n20448, A2 => n19688, B1 => n4890, B2 => 
                           n19699, ZN => n7694);
   U4761 : OAI22_X1 port map( A1 => n20451, A2 => n19688, B1 => n4889, B2 => 
                           n19698, ZN => n7695);
   U4762 : OAI22_X1 port map( A1 => n20454, A2 => n19688, B1 => n4888, B2 => 
                           n19698, ZN => n7696);
   U4763 : OAI22_X1 port map( A1 => n20457, A2 => n19688, B1 => n4887, B2 => 
                           n19698, ZN => n7697);
   U4764 : OAI22_X1 port map( A1 => n20460, A2 => n19688, B1 => n4886, B2 => 
                           n19698, ZN => n7698);
   U4765 : OAI22_X1 port map( A1 => n20463, A2 => n19688, B1 => n4885, B2 => 
                           n19697, ZN => n7699);
   U4766 : OAI22_X1 port map( A1 => n20466, A2 => n19688, B1 => n4884, B2 => 
                           n19697, ZN => n7700);
   U4767 : OAI22_X1 port map( A1 => n20469, A2 => n19688, B1 => n4883, B2 => 
                           n19697, ZN => n7701);
   U4768 : OAI22_X1 port map( A1 => n20472, A2 => n19688, B1 => n4882, B2 => 
                           n19697, ZN => n7702);
   U4769 : OAI22_X1 port map( A1 => n20475, A2 => n19690, B1 => n4881, B2 => 
                           n19696, ZN => n7703);
   U4770 : OAI22_X1 port map( A1 => n20478, A2 => n19689, B1 => n4880, B2 => 
                           n19696, ZN => n7704);
   U4771 : OAI22_X1 port map( A1 => n20481, A2 => n19688, B1 => n4879, B2 => 
                           n19696, ZN => n7705);
   U4772 : OAI22_X1 port map( A1 => n20484, A2 => n19690, B1 => n4878, B2 => 
                           n19696, ZN => n7706);
   U4773 : OAI22_X1 port map( A1 => n20487, A2 => n19689, B1 => n4877, B2 => 
                           n19695, ZN => n7707);
   U4774 : OAI22_X1 port map( A1 => n20490, A2 => n19688, B1 => n4876, B2 => 
                           n19695, ZN => n7708);
   U4775 : OAI22_X1 port map( A1 => n20493, A2 => n19690, B1 => n4875, B2 => 
                           n19695, ZN => n7709);
   U4776 : OAI22_X1 port map( A1 => n20496, A2 => n19689, B1 => n4874, B2 => 
                           n19695, ZN => n7710);
   U4777 : OAI22_X1 port map( A1 => n20499, A2 => n19688, B1 => n4873, B2 => 
                           n19694, ZN => n7711);
   U4778 : OAI22_X1 port map( A1 => n20502, A2 => n19690, B1 => n4872, B2 => 
                           n19694, ZN => n7712);
   U4779 : OAI22_X1 port map( A1 => n20505, A2 => n19689, B1 => n4871, B2 => 
                           n19694, ZN => n7713);
   U4780 : OAI22_X1 port map( A1 => n20508, A2 => n19689, B1 => n4870, B2 => 
                           n19694, ZN => n7714);
   U4781 : OAI22_X1 port map( A1 => n20511, A2 => n19690, B1 => n4869, B2 => 
                           n19693, ZN => n7715);
   U4782 : OAI22_X1 port map( A1 => n20514, A2 => n19689, B1 => n4868, B2 => 
                           n19693, ZN => n7716);
   U4783 : OAI22_X1 port map( A1 => n20517, A2 => n19688, B1 => n4867, B2 => 
                           n19693, ZN => n7717);
   U4784 : OAI22_X1 port map( A1 => n20520, A2 => n19688, B1 => n4866, B2 => 
                           n19693, ZN => n7718);
   U4785 : OAI22_X1 port map( A1 => n20523, A2 => n19690, B1 => n4865, B2 => 
                           n19692, ZN => n7719);
   U4786 : OAI22_X1 port map( A1 => n20526, A2 => n19689, B1 => n4864, B2 => 
                           n19692, ZN => n7720);
   U4787 : OAI22_X1 port map( A1 => n20529, A2 => n19688, B1 => n4863, B2 => 
                           n19692, ZN => n7721);
   U4788 : OAI22_X1 port map( A1 => n20532, A2 => n19690, B1 => n4862, B2 => 
                           n19692, ZN => n7722);
   U4789 : OAI22_X1 port map( A1 => n20535, A2 => n19690, B1 => n4861, B2 => 
                           n19691, ZN => n7723);
   U4790 : OAI22_X1 port map( A1 => n20538, A2 => n19689, B1 => n4860, B2 => 
                           n19691, ZN => n7724);
   U4791 : OAI22_X1 port map( A1 => n20541, A2 => n19688, B1 => n4859, B2 => 
                           n19691, ZN => n7725);
   U4792 : OAI22_X1 port map( A1 => n20572, A2 => n19689, B1 => n4858, B2 => 
                           n19691, ZN => n7726);
   U4793 : OAI22_X1 port map( A1 => n20355, A2 => n19689, B1 => n4921, B2 => 
                           n19706, ZN => n7663);
   U4794 : OAI22_X1 port map( A1 => n20358, A2 => n19688, B1 => n4920, B2 => 
                           n19706, ZN => n7664);
   U4795 : OAI22_X1 port map( A1 => n20361, A2 => n19688, B1 => n4919, B2 => 
                           n19706, ZN => n7665);
   U4796 : OAI22_X1 port map( A1 => n20364, A2 => n19690, B1 => n4918, B2 => 
                           n19706, ZN => n7666);
   U4797 : INV_X1 port map( A => cwp(0), ZN => n11753);
   U4798 : OAI22_X1 port map( A1 => n20369, A2 => n20222, B1 => n3633, B2 => 
                           n20237, ZN => n8883);
   U4799 : OAI22_X1 port map( A1 => n20372, A2 => n20222, B1 => n3632, B2 => 
                           n20237, ZN => n8884);
   U4800 : OAI22_X1 port map( A1 => n20375, A2 => n20222, B1 => n3631, B2 => 
                           n20237, ZN => n8885);
   U4801 : OAI22_X1 port map( A1 => n20378, A2 => n20222, B1 => n3630, B2 => 
                           n20237, ZN => n8886);
   U4802 : OAI22_X1 port map( A1 => n20381, A2 => n20222, B1 => n3629, B2 => 
                           n20236, ZN => n8887);
   U4803 : OAI22_X1 port map( A1 => n20384, A2 => n20222, B1 => n3628, B2 => 
                           n20236, ZN => n8888);
   U4804 : OAI22_X1 port map( A1 => n20387, A2 => n20222, B1 => n3627, B2 => 
                           n20236, ZN => n8889);
   U4805 : OAI22_X1 port map( A1 => n20390, A2 => n20222, B1 => n3626, B2 => 
                           n20236, ZN => n8890);
   U4806 : OAI22_X1 port map( A1 => n20393, A2 => n20222, B1 => n3625, B2 => 
                           n20235, ZN => n8891);
   U4807 : OAI22_X1 port map( A1 => n20396, A2 => n20222, B1 => n3624, B2 => 
                           n20235, ZN => n8892);
   U4808 : OAI22_X1 port map( A1 => n20399, A2 => n20222, B1 => n3623, B2 => 
                           n20235, ZN => n8893);
   U4809 : OAI22_X1 port map( A1 => n20402, A2 => n20222, B1 => n3622, B2 => 
                           n20235, ZN => n8894);
   U4810 : OAI22_X1 port map( A1 => n20405, A2 => n20221, B1 => n3621, B2 => 
                           n20234, ZN => n8895);
   U4811 : OAI22_X1 port map( A1 => n20408, A2 => n20221, B1 => n3620, B2 => 
                           n20234, ZN => n8896);
   U4812 : OAI22_X1 port map( A1 => n20411, A2 => n20221, B1 => n3619, B2 => 
                           n20234, ZN => n8897);
   U4813 : OAI22_X1 port map( A1 => n20414, A2 => n20221, B1 => n3618, B2 => 
                           n20234, ZN => n8898);
   U4814 : OAI22_X1 port map( A1 => n20417, A2 => n20221, B1 => n3617, B2 => 
                           n20233, ZN => n8899);
   U4815 : OAI22_X1 port map( A1 => n20420, A2 => n20221, B1 => n3616, B2 => 
                           n20233, ZN => n8900);
   U4816 : OAI22_X1 port map( A1 => n20423, A2 => n20221, B1 => n3615, B2 => 
                           n20233, ZN => n8901);
   U4817 : OAI22_X1 port map( A1 => n20426, A2 => n20221, B1 => n3614, B2 => 
                           n20233, ZN => n8902);
   U4818 : OAI22_X1 port map( A1 => n20429, A2 => n20221, B1 => n3613, B2 => 
                           n20232, ZN => n8903);
   U4819 : OAI22_X1 port map( A1 => n20432, A2 => n20221, B1 => n3612, B2 => 
                           n20232, ZN => n8904);
   U4820 : OAI22_X1 port map( A1 => n20435, A2 => n20221, B1 => n3611, B2 => 
                           n20232, ZN => n8905);
   U4821 : OAI22_X1 port map( A1 => n20438, A2 => n20221, B1 => n3610, B2 => 
                           n20232, ZN => n8906);
   U4822 : OAI22_X1 port map( A1 => n20441, A2 => n20220, B1 => n3609, B2 => 
                           n20231, ZN => n8907);
   U4823 : OAI22_X1 port map( A1 => n20444, A2 => n20220, B1 => n3608, B2 => 
                           n20231, ZN => n8908);
   U4824 : OAI22_X1 port map( A1 => n20447, A2 => n20220, B1 => n3607, B2 => 
                           n20231, ZN => n8909);
   U4825 : OAI22_X1 port map( A1 => n20450, A2 => n20220, B1 => n3606, B2 => 
                           n20231, ZN => n8910);
   U4826 : OAI22_X1 port map( A1 => n20453, A2 => n20220, B1 => n3605, B2 => 
                           n20230, ZN => n8911);
   U4827 : OAI22_X1 port map( A1 => n20456, A2 => n20220, B1 => n3604, B2 => 
                           n20230, ZN => n8912);
   U4828 : OAI22_X1 port map( A1 => n20459, A2 => n20220, B1 => n3603, B2 => 
                           n20230, ZN => n8913);
   U4829 : OAI22_X1 port map( A1 => n20462, A2 => n20220, B1 => n3602, B2 => 
                           n20230, ZN => n8914);
   U4830 : OAI22_X1 port map( A1 => n20465, A2 => n20220, B1 => n3601, B2 => 
                           n20229, ZN => n8915);
   U4831 : OAI22_X1 port map( A1 => n20468, A2 => n20220, B1 => n3600, B2 => 
                           n20229, ZN => n8916);
   U4832 : OAI22_X1 port map( A1 => n20471, A2 => n20220, B1 => n3599, B2 => 
                           n20229, ZN => n8917);
   U4833 : OAI22_X1 port map( A1 => n20474, A2 => n20220, B1 => n3598, B2 => 
                           n20229, ZN => n8918);
   U4834 : OAI22_X1 port map( A1 => n20477, A2 => n20222, B1 => n3597, B2 => 
                           n20228, ZN => n8919);
   U4835 : OAI22_X1 port map( A1 => n20480, A2 => n20221, B1 => n3596, B2 => 
                           n20228, ZN => n8920);
   U4836 : OAI22_X1 port map( A1 => n20483, A2 => n20220, B1 => n3595, B2 => 
                           n20228, ZN => n8921);
   U4837 : OAI22_X1 port map( A1 => n20486, A2 => n20222, B1 => n3594, B2 => 
                           n20228, ZN => n8922);
   U4838 : OAI22_X1 port map( A1 => n20489, A2 => n20221, B1 => n3593, B2 => 
                           n20227, ZN => n8923);
   U4839 : OAI22_X1 port map( A1 => n20492, A2 => n20220, B1 => n3592, B2 => 
                           n20227, ZN => n8924);
   U4840 : OAI22_X1 port map( A1 => n20495, A2 => n20222, B1 => n3591, B2 => 
                           n20227, ZN => n8925);
   U4841 : OAI22_X1 port map( A1 => n20498, A2 => n20221, B1 => n3590, B2 => 
                           n20227, ZN => n8926);
   U4842 : OAI22_X1 port map( A1 => n20501, A2 => n20220, B1 => n3589, B2 => 
                           n20226, ZN => n8927);
   U4843 : OAI22_X1 port map( A1 => n20504, A2 => n20222, B1 => n3588, B2 => 
                           n20226, ZN => n8928);
   U4844 : OAI22_X1 port map( A1 => n20507, A2 => n20221, B1 => n3587, B2 => 
                           n20226, ZN => n8929);
   U4845 : OAI22_X1 port map( A1 => n20510, A2 => n20221, B1 => n3586, B2 => 
                           n20226, ZN => n8930);
   U4846 : OAI22_X1 port map( A1 => n20513, A2 => n20222, B1 => n3585, B2 => 
                           n20225, ZN => n8931);
   U4847 : OAI22_X1 port map( A1 => n20516, A2 => n20221, B1 => n3584, B2 => 
                           n20225, ZN => n8932);
   U4848 : OAI22_X1 port map( A1 => n20519, A2 => n20220, B1 => n3583, B2 => 
                           n20225, ZN => n8933);
   U4849 : OAI22_X1 port map( A1 => n20522, A2 => n20220, B1 => n3582, B2 => 
                           n20225, ZN => n8934);
   U4850 : OAI22_X1 port map( A1 => n20525, A2 => n20222, B1 => n3581, B2 => 
                           n20224, ZN => n8935);
   U4851 : OAI22_X1 port map( A1 => n20528, A2 => n20221, B1 => n3580, B2 => 
                           n20224, ZN => n8936);
   U4852 : OAI22_X1 port map( A1 => n20531, A2 => n20220, B1 => n3579, B2 => 
                           n20224, ZN => n8937);
   U4853 : OAI22_X1 port map( A1 => n20534, A2 => n20222, B1 => n3578, B2 => 
                           n20224, ZN => n8938);
   U4854 : OAI22_X1 port map( A1 => n20537, A2 => n20222, B1 => n3577, B2 => 
                           n20223, ZN => n8939);
   U4855 : OAI22_X1 port map( A1 => n20540, A2 => n20221, B1 => n3576, B2 => 
                           n20223, ZN => n8940);
   U4856 : OAI22_X1 port map( A1 => n20543, A2 => n20220, B1 => n3575, B2 => 
                           n20223, ZN => n8941);
   U4857 : OAI22_X1 port map( A1 => n20574, A2 => n20221, B1 => n3574, B2 => 
                           n20223, ZN => n8942);
   U4858 : OAI22_X1 port map( A1 => n20357, A2 => n20221, B1 => n3637, B2 => 
                           n20238, ZN => n8879);
   U4859 : OAI22_X1 port map( A1 => n20360, A2 => n20220, B1 => n3636, B2 => 
                           n20238, ZN => n8880);
   U4860 : OAI22_X1 port map( A1 => n20363, A2 => n20220, B1 => n3635, B2 => 
                           n20238, ZN => n8881);
   U4861 : OAI22_X1 port map( A1 => n20366, A2 => n20222, B1 => n3634, B2 => 
                           n20238, ZN => n8882);
   U4862 : OAI22_X1 port map( A1 => n20368, A2 => n20138, B1 => n3832, B2 => 
                           n20153, ZN => n8691);
   U4863 : OAI22_X1 port map( A1 => n20371, A2 => n20138, B1 => n3831, B2 => 
                           n20153, ZN => n8692);
   U4864 : OAI22_X1 port map( A1 => n20374, A2 => n20138, B1 => n3830, B2 => 
                           n20153, ZN => n8693);
   U4865 : OAI22_X1 port map( A1 => n20377, A2 => n20138, B1 => n3829, B2 => 
                           n20153, ZN => n8694);
   U4866 : OAI22_X1 port map( A1 => n20380, A2 => n20138, B1 => n3828, B2 => 
                           n20152, ZN => n8695);
   U4867 : OAI22_X1 port map( A1 => n20383, A2 => n20138, B1 => n3827, B2 => 
                           n20152, ZN => n8696);
   U4868 : OAI22_X1 port map( A1 => n20386, A2 => n20138, B1 => n3826, B2 => 
                           n20152, ZN => n8697);
   U4869 : OAI22_X1 port map( A1 => n20389, A2 => n20138, B1 => n3825, B2 => 
                           n20152, ZN => n8698);
   U4870 : OAI22_X1 port map( A1 => n20392, A2 => n20138, B1 => n3824, B2 => 
                           n20151, ZN => n8699);
   U4871 : OAI22_X1 port map( A1 => n20395, A2 => n20138, B1 => n3823, B2 => 
                           n20151, ZN => n8700);
   U4872 : OAI22_X1 port map( A1 => n20398, A2 => n20138, B1 => n3822, B2 => 
                           n20151, ZN => n8701);
   U4873 : OAI22_X1 port map( A1 => n20401, A2 => n20138, B1 => n3821, B2 => 
                           n20151, ZN => n8702);
   U4874 : OAI22_X1 port map( A1 => n20404, A2 => n20137, B1 => n3820, B2 => 
                           n20150, ZN => n8703);
   U4875 : OAI22_X1 port map( A1 => n20407, A2 => n20137, B1 => n3819, B2 => 
                           n20150, ZN => n8704);
   U4876 : OAI22_X1 port map( A1 => n20410, A2 => n20137, B1 => n3818, B2 => 
                           n20150, ZN => n8705);
   U4877 : OAI22_X1 port map( A1 => n20413, A2 => n20137, B1 => n3817, B2 => 
                           n20150, ZN => n8706);
   U4878 : OAI22_X1 port map( A1 => n20416, A2 => n20137, B1 => n3816, B2 => 
                           n20149, ZN => n8707);
   U4879 : OAI22_X1 port map( A1 => n20419, A2 => n20137, B1 => n3815, B2 => 
                           n20149, ZN => n8708);
   U4880 : OAI22_X1 port map( A1 => n20422, A2 => n20137, B1 => n3814, B2 => 
                           n20149, ZN => n8709);
   U4881 : OAI22_X1 port map( A1 => n20425, A2 => n20137, B1 => n3813, B2 => 
                           n20149, ZN => n8710);
   U4882 : OAI22_X1 port map( A1 => n20428, A2 => n20137, B1 => n3812, B2 => 
                           n20148, ZN => n8711);
   U4883 : OAI22_X1 port map( A1 => n20431, A2 => n20137, B1 => n3811, B2 => 
                           n20148, ZN => n8712);
   U4884 : OAI22_X1 port map( A1 => n20434, A2 => n20137, B1 => n3810, B2 => 
                           n20148, ZN => n8713);
   U4885 : OAI22_X1 port map( A1 => n20437, A2 => n20137, B1 => n3809, B2 => 
                           n20148, ZN => n8714);
   U4886 : OAI22_X1 port map( A1 => n20440, A2 => n20136, B1 => n3808, B2 => 
                           n20147, ZN => n8715);
   U4887 : OAI22_X1 port map( A1 => n20443, A2 => n20136, B1 => n3807, B2 => 
                           n20147, ZN => n8716);
   U4888 : OAI22_X1 port map( A1 => n20446, A2 => n20136, B1 => n3806, B2 => 
                           n20147, ZN => n8717);
   U4889 : OAI22_X1 port map( A1 => n20449, A2 => n20136, B1 => n3805, B2 => 
                           n20147, ZN => n8718);
   U4890 : OAI22_X1 port map( A1 => n20452, A2 => n20136, B1 => n3804, B2 => 
                           n20146, ZN => n8719);
   U4891 : OAI22_X1 port map( A1 => n20455, A2 => n20136, B1 => n3803, B2 => 
                           n20146, ZN => n8720);
   U4892 : OAI22_X1 port map( A1 => n20458, A2 => n20136, B1 => n3802, B2 => 
                           n20146, ZN => n8721);
   U4893 : OAI22_X1 port map( A1 => n20461, A2 => n20136, B1 => n3801, B2 => 
                           n20146, ZN => n8722);
   U4894 : OAI22_X1 port map( A1 => n20464, A2 => n20136, B1 => n3800, B2 => 
                           n20145, ZN => n8723);
   U4895 : OAI22_X1 port map( A1 => n20467, A2 => n20136, B1 => n3799, B2 => 
                           n20145, ZN => n8724);
   U4896 : OAI22_X1 port map( A1 => n20470, A2 => n20136, B1 => n3798, B2 => 
                           n20145, ZN => n8725);
   U4897 : OAI22_X1 port map( A1 => n20473, A2 => n20136, B1 => n3797, B2 => 
                           n20145, ZN => n8726);
   U4898 : OAI22_X1 port map( A1 => n20476, A2 => n20138, B1 => n3796, B2 => 
                           n20144, ZN => n8727);
   U4899 : OAI22_X1 port map( A1 => n20479, A2 => n20137, B1 => n3795, B2 => 
                           n20144, ZN => n8728);
   U4900 : OAI22_X1 port map( A1 => n20482, A2 => n20136, B1 => n3794, B2 => 
                           n20144, ZN => n8729);
   U4901 : OAI22_X1 port map( A1 => n20485, A2 => n20138, B1 => n3793, B2 => 
                           n20144, ZN => n8730);
   U4902 : OAI22_X1 port map( A1 => n20488, A2 => n20137, B1 => n3792, B2 => 
                           n20143, ZN => n8731);
   U4903 : OAI22_X1 port map( A1 => n20491, A2 => n20136, B1 => n3791, B2 => 
                           n20143, ZN => n8732);
   U4904 : OAI22_X1 port map( A1 => n20494, A2 => n20138, B1 => n3790, B2 => 
                           n20143, ZN => n8733);
   U4905 : OAI22_X1 port map( A1 => n20497, A2 => n20137, B1 => n3789, B2 => 
                           n20143, ZN => n8734);
   U4906 : OAI22_X1 port map( A1 => n20500, A2 => n20136, B1 => n3788, B2 => 
                           n20142, ZN => n8735);
   U4907 : OAI22_X1 port map( A1 => n20503, A2 => n20138, B1 => n3787, B2 => 
                           n20142, ZN => n8736);
   U4908 : OAI22_X1 port map( A1 => n20506, A2 => n20137, B1 => n3786, B2 => 
                           n20142, ZN => n8737);
   U4909 : OAI22_X1 port map( A1 => n20509, A2 => n20137, B1 => n3785, B2 => 
                           n20142, ZN => n8738);
   U4910 : OAI22_X1 port map( A1 => n20512, A2 => n20138, B1 => n3784, B2 => 
                           n20141, ZN => n8739);
   U4911 : OAI22_X1 port map( A1 => n20515, A2 => n20137, B1 => n3783, B2 => 
                           n20141, ZN => n8740);
   U4912 : OAI22_X1 port map( A1 => n20518, A2 => n20136, B1 => n3782, B2 => 
                           n20141, ZN => n8741);
   U4913 : OAI22_X1 port map( A1 => n20521, A2 => n20136, B1 => n3781, B2 => 
                           n20141, ZN => n8742);
   U4914 : OAI22_X1 port map( A1 => n20524, A2 => n20138, B1 => n3780, B2 => 
                           n20140, ZN => n8743);
   U4915 : OAI22_X1 port map( A1 => n20527, A2 => n20137, B1 => n3779, B2 => 
                           n20140, ZN => n8744);
   U4916 : OAI22_X1 port map( A1 => n20530, A2 => n20136, B1 => n3778, B2 => 
                           n20140, ZN => n8745);
   U4917 : OAI22_X1 port map( A1 => n20533, A2 => n20138, B1 => n3777, B2 => 
                           n20140, ZN => n8746);
   U4918 : OAI22_X1 port map( A1 => n20536, A2 => n20138, B1 => n3776, B2 => 
                           n20139, ZN => n8747);
   U4919 : OAI22_X1 port map( A1 => n20539, A2 => n20137, B1 => n3775, B2 => 
                           n20139, ZN => n8748);
   U4920 : OAI22_X1 port map( A1 => n20542, A2 => n20136, B1 => n3774, B2 => 
                           n20139, ZN => n8749);
   U4921 : OAI22_X1 port map( A1 => n20573, A2 => n20137, B1 => n3773, B2 => 
                           n20139, ZN => n8750);
   U4922 : OAI22_X1 port map( A1 => n20356, A2 => n20137, B1 => n3836, B2 => 
                           n20154, ZN => n8687);
   U4923 : OAI22_X1 port map( A1 => n20359, A2 => n20136, B1 => n3835, B2 => 
                           n20154, ZN => n8688);
   U4924 : OAI22_X1 port map( A1 => n20362, A2 => n20136, B1 => n3834, B2 => 
                           n20154, ZN => n8689);
   U4925 : OAI22_X1 port map( A1 => n20365, A2 => n20138, B1 => n3833, B2 => 
                           n20154, ZN => n8690);
   U4926 : OAI22_X1 port map( A1 => n20368, A2 => n19858, B1 => n4507, B2 => 
                           n19873, ZN => n8051);
   U4927 : OAI22_X1 port map( A1 => n20371, A2 => n19858, B1 => n4506, B2 => 
                           n19873, ZN => n8052);
   U4928 : OAI22_X1 port map( A1 => n20374, A2 => n19858, B1 => n4505, B2 => 
                           n19873, ZN => n8053);
   U4929 : OAI22_X1 port map( A1 => n20377, A2 => n19858, B1 => n4504, B2 => 
                           n19873, ZN => n8054);
   U4930 : OAI22_X1 port map( A1 => n20380, A2 => n19858, B1 => n4503, B2 => 
                           n19872, ZN => n8055);
   U4931 : OAI22_X1 port map( A1 => n20383, A2 => n19858, B1 => n4502, B2 => 
                           n19872, ZN => n8056);
   U4932 : OAI22_X1 port map( A1 => n20386, A2 => n19858, B1 => n4501, B2 => 
                           n19872, ZN => n8057);
   U4933 : OAI22_X1 port map( A1 => n20389, A2 => n19858, B1 => n4500, B2 => 
                           n19872, ZN => n8058);
   U4934 : OAI22_X1 port map( A1 => n20392, A2 => n19858, B1 => n4499, B2 => 
                           n19871, ZN => n8059);
   U4935 : OAI22_X1 port map( A1 => n20395, A2 => n19858, B1 => n4498, B2 => 
                           n19871, ZN => n8060);
   U4936 : OAI22_X1 port map( A1 => n20398, A2 => n19858, B1 => n4497, B2 => 
                           n19871, ZN => n8061);
   U4937 : OAI22_X1 port map( A1 => n20401, A2 => n19858, B1 => n4496, B2 => 
                           n19871, ZN => n8062);
   U4938 : OAI22_X1 port map( A1 => n20404, A2 => n19857, B1 => n4495, B2 => 
                           n19870, ZN => n8063);
   U4939 : OAI22_X1 port map( A1 => n20407, A2 => n19857, B1 => n4494, B2 => 
                           n19870, ZN => n8064);
   U4940 : OAI22_X1 port map( A1 => n20410, A2 => n19857, B1 => n4493, B2 => 
                           n19870, ZN => n8065);
   U4941 : OAI22_X1 port map( A1 => n20413, A2 => n19857, B1 => n4492, B2 => 
                           n19870, ZN => n8066);
   U4942 : OAI22_X1 port map( A1 => n20416, A2 => n19857, B1 => n4491, B2 => 
                           n19869, ZN => n8067);
   U4943 : OAI22_X1 port map( A1 => n20419, A2 => n19857, B1 => n4490, B2 => 
                           n19869, ZN => n8068);
   U4944 : OAI22_X1 port map( A1 => n20422, A2 => n19857, B1 => n4489, B2 => 
                           n19869, ZN => n8069);
   U4945 : OAI22_X1 port map( A1 => n20425, A2 => n19857, B1 => n4488, B2 => 
                           n19869, ZN => n8070);
   U4946 : OAI22_X1 port map( A1 => n20428, A2 => n19857, B1 => n4487, B2 => 
                           n19868, ZN => n8071);
   U4947 : OAI22_X1 port map( A1 => n20431, A2 => n19857, B1 => n4486, B2 => 
                           n19868, ZN => n8072);
   U4948 : OAI22_X1 port map( A1 => n20434, A2 => n19857, B1 => n4485, B2 => 
                           n19868, ZN => n8073);
   U4949 : OAI22_X1 port map( A1 => n20437, A2 => n19857, B1 => n4484, B2 => 
                           n19868, ZN => n8074);
   U4950 : OAI22_X1 port map( A1 => n20440, A2 => n19856, B1 => n4483, B2 => 
                           n19867, ZN => n8075);
   U4951 : OAI22_X1 port map( A1 => n20443, A2 => n19856, B1 => n4482, B2 => 
                           n19867, ZN => n8076);
   U4952 : OAI22_X1 port map( A1 => n20446, A2 => n19856, B1 => n4481, B2 => 
                           n19867, ZN => n8077);
   U4953 : OAI22_X1 port map( A1 => n20449, A2 => n19856, B1 => n4480, B2 => 
                           n19867, ZN => n8078);
   U4954 : OAI22_X1 port map( A1 => n20452, A2 => n19856, B1 => n4479, B2 => 
                           n19866, ZN => n8079);
   U4955 : OAI22_X1 port map( A1 => n20455, A2 => n19856, B1 => n4478, B2 => 
                           n19866, ZN => n8080);
   U4956 : OAI22_X1 port map( A1 => n20458, A2 => n19856, B1 => n4477, B2 => 
                           n19866, ZN => n8081);
   U4957 : OAI22_X1 port map( A1 => n20461, A2 => n19856, B1 => n4476, B2 => 
                           n19866, ZN => n8082);
   U4958 : OAI22_X1 port map( A1 => n20464, A2 => n19856, B1 => n4475, B2 => 
                           n19865, ZN => n8083);
   U4959 : OAI22_X1 port map( A1 => n20467, A2 => n19856, B1 => n4474, B2 => 
                           n19865, ZN => n8084);
   U4960 : OAI22_X1 port map( A1 => n20470, A2 => n19856, B1 => n4473, B2 => 
                           n19865, ZN => n8085);
   U4961 : OAI22_X1 port map( A1 => n20473, A2 => n19856, B1 => n4472, B2 => 
                           n19865, ZN => n8086);
   U4962 : OAI22_X1 port map( A1 => n20476, A2 => n19858, B1 => n4471, B2 => 
                           n19864, ZN => n8087);
   U4963 : OAI22_X1 port map( A1 => n20479, A2 => n19857, B1 => n4470, B2 => 
                           n19864, ZN => n8088);
   U4964 : OAI22_X1 port map( A1 => n20482, A2 => n19856, B1 => n4469, B2 => 
                           n19864, ZN => n8089);
   U4965 : OAI22_X1 port map( A1 => n20485, A2 => n19858, B1 => n4468, B2 => 
                           n19864, ZN => n8090);
   U4966 : OAI22_X1 port map( A1 => n20488, A2 => n19857, B1 => n4467, B2 => 
                           n19863, ZN => n8091);
   U4967 : OAI22_X1 port map( A1 => n20491, A2 => n19856, B1 => n4466, B2 => 
                           n19863, ZN => n8092);
   U4968 : OAI22_X1 port map( A1 => n20494, A2 => n19858, B1 => n4465, B2 => 
                           n19863, ZN => n8093);
   U4969 : OAI22_X1 port map( A1 => n20497, A2 => n19857, B1 => n4464, B2 => 
                           n19863, ZN => n8094);
   U4970 : OAI22_X1 port map( A1 => n20500, A2 => n19856, B1 => n4463, B2 => 
                           n19862, ZN => n8095);
   U4971 : OAI22_X1 port map( A1 => n20503, A2 => n19858, B1 => n4462, B2 => 
                           n19862, ZN => n8096);
   U4972 : OAI22_X1 port map( A1 => n20506, A2 => n19857, B1 => n4461, B2 => 
                           n19862, ZN => n8097);
   U4973 : OAI22_X1 port map( A1 => n20509, A2 => n19857, B1 => n4460, B2 => 
                           n19862, ZN => n8098);
   U4974 : OAI22_X1 port map( A1 => n20512, A2 => n19858, B1 => n4459, B2 => 
                           n19861, ZN => n8099);
   U4975 : OAI22_X1 port map( A1 => n20515, A2 => n19857, B1 => n4458, B2 => 
                           n19861, ZN => n8100);
   U4976 : OAI22_X1 port map( A1 => n20518, A2 => n19856, B1 => n4457, B2 => 
                           n19861, ZN => n8101);
   U4977 : OAI22_X1 port map( A1 => n20521, A2 => n19856, B1 => n4456, B2 => 
                           n19861, ZN => n8102);
   U4978 : OAI22_X1 port map( A1 => n20524, A2 => n19858, B1 => n4455, B2 => 
                           n19860, ZN => n8103);
   U4979 : OAI22_X1 port map( A1 => n20527, A2 => n19857, B1 => n4454, B2 => 
                           n19860, ZN => n8104);
   U4980 : OAI22_X1 port map( A1 => n20530, A2 => n19856, B1 => n4453, B2 => 
                           n19860, ZN => n8105);
   U4981 : OAI22_X1 port map( A1 => n20533, A2 => n19858, B1 => n4452, B2 => 
                           n19860, ZN => n8106);
   U4982 : OAI22_X1 port map( A1 => n20536, A2 => n19858, B1 => n4451, B2 => 
                           n19859, ZN => n8107);
   U4983 : OAI22_X1 port map( A1 => n20539, A2 => n19857, B1 => n4450, B2 => 
                           n19859, ZN => n8108);
   U4984 : OAI22_X1 port map( A1 => n20542, A2 => n19856, B1 => n4449, B2 => 
                           n19859, ZN => n8109);
   U4985 : OAI22_X1 port map( A1 => n20573, A2 => n19857, B1 => n4448, B2 => 
                           n19859, ZN => n8110);
   U4986 : OAI22_X1 port map( A1 => n20369, A2 => n20250, B1 => n3565, B2 => 
                           n20265, ZN => n8947);
   U4987 : OAI22_X1 port map( A1 => n20372, A2 => n20250, B1 => n3564, B2 => 
                           n20265, ZN => n8948);
   U4988 : OAI22_X1 port map( A1 => n20375, A2 => n20250, B1 => n3563, B2 => 
                           n20265, ZN => n8949);
   U4989 : OAI22_X1 port map( A1 => n20378, A2 => n20250, B1 => n3562, B2 => 
                           n20265, ZN => n8950);
   U4990 : OAI22_X1 port map( A1 => n20381, A2 => n20250, B1 => n3561, B2 => 
                           n20264, ZN => n8951);
   U4991 : OAI22_X1 port map( A1 => n20384, A2 => n20250, B1 => n3560, B2 => 
                           n20264, ZN => n8952);
   U4992 : OAI22_X1 port map( A1 => n20387, A2 => n20250, B1 => n3559, B2 => 
                           n20264, ZN => n8953);
   U4993 : OAI22_X1 port map( A1 => n20390, A2 => n20250, B1 => n3558, B2 => 
                           n20264, ZN => n8954);
   U4994 : OAI22_X1 port map( A1 => n20393, A2 => n20250, B1 => n3557, B2 => 
                           n20263, ZN => n8955);
   U4995 : OAI22_X1 port map( A1 => n20396, A2 => n20250, B1 => n3556, B2 => 
                           n20263, ZN => n8956);
   U4996 : OAI22_X1 port map( A1 => n20399, A2 => n20250, B1 => n3555, B2 => 
                           n20263, ZN => n8957);
   U4997 : OAI22_X1 port map( A1 => n20402, A2 => n20250, B1 => n3554, B2 => 
                           n20263, ZN => n8958);
   U4998 : OAI22_X1 port map( A1 => n20405, A2 => n20249, B1 => n3553, B2 => 
                           n20262, ZN => n8959);
   U4999 : OAI22_X1 port map( A1 => n20408, A2 => n20249, B1 => n3552, B2 => 
                           n20262, ZN => n8960);
   U5000 : OAI22_X1 port map( A1 => n20411, A2 => n20249, B1 => n3551, B2 => 
                           n20262, ZN => n8961);
   U5001 : OAI22_X1 port map( A1 => n20414, A2 => n20249, B1 => n3550, B2 => 
                           n20262, ZN => n8962);
   U5002 : OAI22_X1 port map( A1 => n20417, A2 => n20249, B1 => n3549, B2 => 
                           n20261, ZN => n8963);
   U5003 : OAI22_X1 port map( A1 => n20420, A2 => n20249, B1 => n3548, B2 => 
                           n20261, ZN => n8964);
   U5004 : OAI22_X1 port map( A1 => n20423, A2 => n20249, B1 => n3547, B2 => 
                           n20261, ZN => n8965);
   U5005 : OAI22_X1 port map( A1 => n20426, A2 => n20249, B1 => n3546, B2 => 
                           n20261, ZN => n8966);
   U5006 : OAI22_X1 port map( A1 => n20429, A2 => n20249, B1 => n3545, B2 => 
                           n20260, ZN => n8967);
   U5007 : OAI22_X1 port map( A1 => n20432, A2 => n20249, B1 => n3544, B2 => 
                           n20260, ZN => n8968);
   U5008 : OAI22_X1 port map( A1 => n20435, A2 => n20249, B1 => n3543, B2 => 
                           n20260, ZN => n8969);
   U5009 : OAI22_X1 port map( A1 => n20438, A2 => n20249, B1 => n3542, B2 => 
                           n20260, ZN => n8970);
   U5010 : OAI22_X1 port map( A1 => n20441, A2 => n20248, B1 => n3541, B2 => 
                           n20259, ZN => n8971);
   U5011 : OAI22_X1 port map( A1 => n20444, A2 => n20248, B1 => n3540, B2 => 
                           n20259, ZN => n8972);
   U5012 : OAI22_X1 port map( A1 => n20447, A2 => n20248, B1 => n3539, B2 => 
                           n20259, ZN => n8973);
   U5013 : OAI22_X1 port map( A1 => n20450, A2 => n20248, B1 => n3538, B2 => 
                           n20259, ZN => n8974);
   U5014 : OAI22_X1 port map( A1 => n20453, A2 => n20248, B1 => n3537, B2 => 
                           n20258, ZN => n8975);
   U5015 : OAI22_X1 port map( A1 => n20456, A2 => n20248, B1 => n3536, B2 => 
                           n20258, ZN => n8976);
   U5016 : OAI22_X1 port map( A1 => n20459, A2 => n20248, B1 => n3535, B2 => 
                           n20258, ZN => n8977);
   U5017 : OAI22_X1 port map( A1 => n20462, A2 => n20248, B1 => n3534, B2 => 
                           n20258, ZN => n8978);
   U5018 : OAI22_X1 port map( A1 => n20465, A2 => n20248, B1 => n3533, B2 => 
                           n20257, ZN => n8979);
   U5019 : OAI22_X1 port map( A1 => n20468, A2 => n20248, B1 => n3532, B2 => 
                           n20257, ZN => n8980);
   U5020 : OAI22_X1 port map( A1 => n20471, A2 => n20248, B1 => n3531, B2 => 
                           n20257, ZN => n8981);
   U5021 : OAI22_X1 port map( A1 => n20474, A2 => n20248, B1 => n3530, B2 => 
                           n20257, ZN => n8982);
   U5022 : OAI22_X1 port map( A1 => n20477, A2 => n20250, B1 => n3529, B2 => 
                           n20256, ZN => n8983);
   U5023 : OAI22_X1 port map( A1 => n20480, A2 => n20249, B1 => n3528, B2 => 
                           n20256, ZN => n8984);
   U5024 : OAI22_X1 port map( A1 => n20483, A2 => n20248, B1 => n3527, B2 => 
                           n20256, ZN => n8985);
   U5025 : OAI22_X1 port map( A1 => n20486, A2 => n20250, B1 => n3526, B2 => 
                           n20256, ZN => n8986);
   U5026 : OAI22_X1 port map( A1 => n20489, A2 => n20249, B1 => n3525, B2 => 
                           n20255, ZN => n8987);
   U5027 : OAI22_X1 port map( A1 => n20492, A2 => n20248, B1 => n3524, B2 => 
                           n20255, ZN => n8988);
   U5028 : OAI22_X1 port map( A1 => n20495, A2 => n20250, B1 => n3523, B2 => 
                           n20255, ZN => n8989);
   U5029 : OAI22_X1 port map( A1 => n20498, A2 => n20249, B1 => n3522, B2 => 
                           n20255, ZN => n8990);
   U5030 : OAI22_X1 port map( A1 => n20501, A2 => n20248, B1 => n3521, B2 => 
                           n20254, ZN => n8991);
   U5031 : OAI22_X1 port map( A1 => n20504, A2 => n20250, B1 => n3520, B2 => 
                           n20254, ZN => n8992);
   U5032 : OAI22_X1 port map( A1 => n20507, A2 => n20249, B1 => n3519, B2 => 
                           n20254, ZN => n8993);
   U5033 : OAI22_X1 port map( A1 => n20510, A2 => n20249, B1 => n3518, B2 => 
                           n20254, ZN => n8994);
   U5034 : OAI22_X1 port map( A1 => n20513, A2 => n20250, B1 => n3517, B2 => 
                           n20253, ZN => n8995);
   U5035 : OAI22_X1 port map( A1 => n20516, A2 => n20249, B1 => n3516, B2 => 
                           n20253, ZN => n8996);
   U5036 : OAI22_X1 port map( A1 => n20519, A2 => n20248, B1 => n3515, B2 => 
                           n20253, ZN => n8997);
   U5037 : OAI22_X1 port map( A1 => n20522, A2 => n20248, B1 => n3514, B2 => 
                           n20253, ZN => n8998);
   U5038 : OAI22_X1 port map( A1 => n20525, A2 => n20250, B1 => n3513, B2 => 
                           n20252, ZN => n8999);
   U5039 : OAI22_X1 port map( A1 => n20528, A2 => n20249, B1 => n3512, B2 => 
                           n20252, ZN => n9000);
   U5040 : OAI22_X1 port map( A1 => n20531, A2 => n20248, B1 => n3511, B2 => 
                           n20252, ZN => n9001);
   U5041 : OAI22_X1 port map( A1 => n20534, A2 => n20250, B1 => n3510, B2 => 
                           n20252, ZN => n9002);
   U5042 : OAI22_X1 port map( A1 => n20537, A2 => n20250, B1 => n3509, B2 => 
                           n20251, ZN => n9003);
   U5043 : OAI22_X1 port map( A1 => n20540, A2 => n20249, B1 => n3508, B2 => 
                           n20251, ZN => n9004);
   U5044 : OAI22_X1 port map( A1 => n20543, A2 => n20248, B1 => n3507, B2 => 
                           n20251, ZN => n9005);
   U5045 : OAI22_X1 port map( A1 => n20574, A2 => n20249, B1 => n3506, B2 => 
                           n20251, ZN => n9006);
   U5046 : OAI22_X1 port map( A1 => n20356, A2 => n19857, B1 => n4511, B2 => 
                           n19874, ZN => n8047);
   U5047 : OAI22_X1 port map( A1 => n20359, A2 => n19856, B1 => n4510, B2 => 
                           n19874, ZN => n8048);
   U5048 : OAI22_X1 port map( A1 => n20362, A2 => n19856, B1 => n4509, B2 => 
                           n19874, ZN => n8049);
   U5049 : OAI22_X1 port map( A1 => n20365, A2 => n19858, B1 => n4508, B2 => 
                           n19874, ZN => n8050);
   U5050 : OAI22_X1 port map( A1 => n20357, A2 => n20249, B1 => n3569, B2 => 
                           n20266, ZN => n8943);
   U5051 : OAI22_X1 port map( A1 => n20360, A2 => n20248, B1 => n3568, B2 => 
                           n20266, ZN => n8944);
   U5052 : OAI22_X1 port map( A1 => n20363, A2 => n20248, B1 => n3567, B2 => 
                           n20266, ZN => n8945);
   U5053 : OAI22_X1 port map( A1 => n20366, A2 => n20250, B1 => n3566, B2 => 
                           n20266, ZN => n8946);
   U5054 : OAI22_X1 port map( A1 => n20367, A2 => n19774, B1 => n4713, B2 => 
                           n19789, ZN => n7859);
   U5055 : OAI22_X1 port map( A1 => n20370, A2 => n19774, B1 => n4712, B2 => 
                           n19789, ZN => n7860);
   U5056 : OAI22_X1 port map( A1 => n20373, A2 => n19774, B1 => n4711, B2 => 
                           n19789, ZN => n7861);
   U5057 : OAI22_X1 port map( A1 => n20376, A2 => n19774, B1 => n4710, B2 => 
                           n19789, ZN => n7862);
   U5058 : OAI22_X1 port map( A1 => n20379, A2 => n19774, B1 => n4709, B2 => 
                           n19788, ZN => n7863);
   U5059 : OAI22_X1 port map( A1 => n20382, A2 => n19774, B1 => n4708, B2 => 
                           n19788, ZN => n7864);
   U5060 : OAI22_X1 port map( A1 => n20385, A2 => n19774, B1 => n4707, B2 => 
                           n19788, ZN => n7865);
   U5061 : OAI22_X1 port map( A1 => n20388, A2 => n19774, B1 => n4706, B2 => 
                           n19788, ZN => n7866);
   U5062 : OAI22_X1 port map( A1 => n20391, A2 => n19774, B1 => n4705, B2 => 
                           n19787, ZN => n7867);
   U5063 : OAI22_X1 port map( A1 => n20394, A2 => n19774, B1 => n4704, B2 => 
                           n19787, ZN => n7868);
   U5064 : OAI22_X1 port map( A1 => n20397, A2 => n19774, B1 => n4703, B2 => 
                           n19787, ZN => n7869);
   U5065 : OAI22_X1 port map( A1 => n20400, A2 => n19774, B1 => n4702, B2 => 
                           n19787, ZN => n7870);
   U5066 : OAI22_X1 port map( A1 => n20403, A2 => n19773, B1 => n4701, B2 => 
                           n19786, ZN => n7871);
   U5067 : OAI22_X1 port map( A1 => n20406, A2 => n19773, B1 => n4700, B2 => 
                           n19786, ZN => n7872);
   U5068 : OAI22_X1 port map( A1 => n20409, A2 => n19773, B1 => n4699, B2 => 
                           n19786, ZN => n7873);
   U5069 : OAI22_X1 port map( A1 => n20412, A2 => n19773, B1 => n4698, B2 => 
                           n19786, ZN => n7874);
   U5070 : OAI22_X1 port map( A1 => n20415, A2 => n19773, B1 => n4697, B2 => 
                           n19785, ZN => n7875);
   U5071 : OAI22_X1 port map( A1 => n20418, A2 => n19773, B1 => n4696, B2 => 
                           n19785, ZN => n7876);
   U5072 : OAI22_X1 port map( A1 => n20421, A2 => n19773, B1 => n4695, B2 => 
                           n19785, ZN => n7877);
   U5073 : OAI22_X1 port map( A1 => n20424, A2 => n19773, B1 => n4694, B2 => 
                           n19785, ZN => n7878);
   U5074 : OAI22_X1 port map( A1 => n20427, A2 => n19773, B1 => n4693, B2 => 
                           n19784, ZN => n7879);
   U5075 : OAI22_X1 port map( A1 => n20430, A2 => n19773, B1 => n4692, B2 => 
                           n19784, ZN => n7880);
   U5076 : OAI22_X1 port map( A1 => n20433, A2 => n19773, B1 => n4691, B2 => 
                           n19784, ZN => n7881);
   U5077 : OAI22_X1 port map( A1 => n20436, A2 => n19773, B1 => n4690, B2 => 
                           n19784, ZN => n7882);
   U5078 : OAI22_X1 port map( A1 => n20439, A2 => n19772, B1 => n4689, B2 => 
                           n19783, ZN => n7883);
   U5079 : OAI22_X1 port map( A1 => n20442, A2 => n19772, B1 => n4688, B2 => 
                           n19783, ZN => n7884);
   U5080 : OAI22_X1 port map( A1 => n20445, A2 => n19772, B1 => n4687, B2 => 
                           n19783, ZN => n7885);
   U5081 : OAI22_X1 port map( A1 => n20448, A2 => n19772, B1 => n4686, B2 => 
                           n19783, ZN => n7886);
   U5082 : OAI22_X1 port map( A1 => n20451, A2 => n19772, B1 => n4685, B2 => 
                           n19782, ZN => n7887);
   U5083 : OAI22_X1 port map( A1 => n20454, A2 => n19772, B1 => n4684, B2 => 
                           n19782, ZN => n7888);
   U5084 : OAI22_X1 port map( A1 => n20457, A2 => n19772, B1 => n4683, B2 => 
                           n19782, ZN => n7889);
   U5085 : OAI22_X1 port map( A1 => n20460, A2 => n19772, B1 => n4682, B2 => 
                           n19782, ZN => n7890);
   U5086 : OAI22_X1 port map( A1 => n20463, A2 => n19772, B1 => n4681, B2 => 
                           n19781, ZN => n7891);
   U5087 : OAI22_X1 port map( A1 => n20466, A2 => n19772, B1 => n4680, B2 => 
                           n19781, ZN => n7892);
   U5088 : OAI22_X1 port map( A1 => n20469, A2 => n19772, B1 => n4679, B2 => 
                           n19781, ZN => n7893);
   U5089 : OAI22_X1 port map( A1 => n20472, A2 => n19772, B1 => n4678, B2 => 
                           n19781, ZN => n7894);
   U5090 : OAI22_X1 port map( A1 => n20475, A2 => n19774, B1 => n4677, B2 => 
                           n19780, ZN => n7895);
   U5091 : OAI22_X1 port map( A1 => n20478, A2 => n19773, B1 => n4676, B2 => 
                           n19780, ZN => n7896);
   U5092 : OAI22_X1 port map( A1 => n20481, A2 => n19772, B1 => n4675, B2 => 
                           n19780, ZN => n7897);
   U5093 : OAI22_X1 port map( A1 => n20484, A2 => n19774, B1 => n4674, B2 => 
                           n19780, ZN => n7898);
   U5094 : OAI22_X1 port map( A1 => n20487, A2 => n19773, B1 => n4673, B2 => 
                           n19779, ZN => n7899);
   U5095 : OAI22_X1 port map( A1 => n20490, A2 => n19772, B1 => n4672, B2 => 
                           n19779, ZN => n7900);
   U5096 : OAI22_X1 port map( A1 => n20493, A2 => n19774, B1 => n4671, B2 => 
                           n19779, ZN => n7901);
   U5097 : OAI22_X1 port map( A1 => n20496, A2 => n19773, B1 => n4670, B2 => 
                           n19779, ZN => n7902);
   U5098 : OAI22_X1 port map( A1 => n20499, A2 => n19772, B1 => n4669, B2 => 
                           n19778, ZN => n7903);
   U5099 : OAI22_X1 port map( A1 => n20502, A2 => n19774, B1 => n4668, B2 => 
                           n19778, ZN => n7904);
   U5100 : OAI22_X1 port map( A1 => n20505, A2 => n19773, B1 => n4667, B2 => 
                           n19778, ZN => n7905);
   U5101 : OAI22_X1 port map( A1 => n20508, A2 => n19773, B1 => n4666, B2 => 
                           n19778, ZN => n7906);
   U5102 : OAI22_X1 port map( A1 => n20511, A2 => n19774, B1 => n4665, B2 => 
                           n19777, ZN => n7907);
   U5103 : OAI22_X1 port map( A1 => n20514, A2 => n19773, B1 => n4664, B2 => 
                           n19777, ZN => n7908);
   U5104 : OAI22_X1 port map( A1 => n20517, A2 => n19772, B1 => n4663, B2 => 
                           n19777, ZN => n7909);
   U5105 : OAI22_X1 port map( A1 => n20520, A2 => n19772, B1 => n4662, B2 => 
                           n19777, ZN => n7910);
   U5106 : OAI22_X1 port map( A1 => n20523, A2 => n19774, B1 => n4661, B2 => 
                           n19776, ZN => n7911);
   U5107 : OAI22_X1 port map( A1 => n20526, A2 => n19773, B1 => n4660, B2 => 
                           n19776, ZN => n7912);
   U5108 : OAI22_X1 port map( A1 => n20529, A2 => n19772, B1 => n4659, B2 => 
                           n19776, ZN => n7913);
   U5109 : OAI22_X1 port map( A1 => n20532, A2 => n19774, B1 => n4658, B2 => 
                           n19776, ZN => n7914);
   U5110 : OAI22_X1 port map( A1 => n20535, A2 => n19774, B1 => n4657, B2 => 
                           n19775, ZN => n7915);
   U5111 : OAI22_X1 port map( A1 => n20538, A2 => n19773, B1 => n4656, B2 => 
                           n19775, ZN => n7916);
   U5112 : OAI22_X1 port map( A1 => n20541, A2 => n19772, B1 => n4655, B2 => 
                           n19775, ZN => n7917);
   U5113 : OAI22_X1 port map( A1 => n20572, A2 => n19773, B1 => n4654, B2 => 
                           n19775, ZN => n7918);
   U5114 : OAI22_X1 port map( A1 => n20355, A2 => n19773, B1 => n4717, B2 => 
                           n19790, ZN => n7855);
   U5115 : OAI22_X1 port map( A1 => n20358, A2 => n19772, B1 => n4716, B2 => 
                           n19790, ZN => n7856);
   U5116 : OAI22_X1 port map( A1 => n20361, A2 => n19772, B1 => n4715, B2 => 
                           n19790, ZN => n7857);
   U5117 : OAI22_X1 port map( A1 => n20364, A2 => n19774, B1 => n4714, B2 => 
                           n19790, ZN => n7858);
   U5118 : OAI22_X1 port map( A1 => n20368, A2 => n19970, B1 => n4238, B2 => 
                           n19985, ZN => n8307);
   U5119 : OAI22_X1 port map( A1 => n20371, A2 => n19970, B1 => n4237, B2 => 
                           n19985, ZN => n8308);
   U5120 : OAI22_X1 port map( A1 => n20374, A2 => n19970, B1 => n4236, B2 => 
                           n19985, ZN => n8309);
   U5121 : OAI22_X1 port map( A1 => n20377, A2 => n19970, B1 => n4235, B2 => 
                           n19985, ZN => n8310);
   U5122 : OAI22_X1 port map( A1 => n20380, A2 => n19970, B1 => n4234, B2 => 
                           n19984, ZN => n8311);
   U5123 : OAI22_X1 port map( A1 => n20383, A2 => n19970, B1 => n4233, B2 => 
                           n19984, ZN => n8312);
   U5124 : OAI22_X1 port map( A1 => n20386, A2 => n19970, B1 => n4232, B2 => 
                           n19984, ZN => n8313);
   U5125 : OAI22_X1 port map( A1 => n20389, A2 => n19970, B1 => n4231, B2 => 
                           n19984, ZN => n8314);
   U5126 : OAI22_X1 port map( A1 => n20392, A2 => n19970, B1 => n4230, B2 => 
                           n19983, ZN => n8315);
   U5127 : OAI22_X1 port map( A1 => n20395, A2 => n19970, B1 => n4229, B2 => 
                           n19983, ZN => n8316);
   U5128 : OAI22_X1 port map( A1 => n20398, A2 => n19970, B1 => n4228, B2 => 
                           n19983, ZN => n8317);
   U5129 : OAI22_X1 port map( A1 => n20401, A2 => n19970, B1 => n4227, B2 => 
                           n19983, ZN => n8318);
   U5130 : OAI22_X1 port map( A1 => n20404, A2 => n19969, B1 => n4226, B2 => 
                           n19982, ZN => n8319);
   U5131 : OAI22_X1 port map( A1 => n20407, A2 => n19969, B1 => n4225, B2 => 
                           n19982, ZN => n8320);
   U5132 : OAI22_X1 port map( A1 => n20410, A2 => n19969, B1 => n4224, B2 => 
                           n19982, ZN => n8321);
   U5133 : OAI22_X1 port map( A1 => n20413, A2 => n19969, B1 => n4223, B2 => 
                           n19982, ZN => n8322);
   U5134 : OAI22_X1 port map( A1 => n20416, A2 => n19969, B1 => n4222, B2 => 
                           n19981, ZN => n8323);
   U5135 : OAI22_X1 port map( A1 => n20419, A2 => n19969, B1 => n4221, B2 => 
                           n19981, ZN => n8324);
   U5136 : OAI22_X1 port map( A1 => n20422, A2 => n19969, B1 => n4220, B2 => 
                           n19981, ZN => n8325);
   U5137 : OAI22_X1 port map( A1 => n20425, A2 => n19969, B1 => n4219, B2 => 
                           n19981, ZN => n8326);
   U5138 : OAI22_X1 port map( A1 => n20428, A2 => n19969, B1 => n4218, B2 => 
                           n19980, ZN => n8327);
   U5139 : OAI22_X1 port map( A1 => n20431, A2 => n19969, B1 => n4217, B2 => 
                           n19980, ZN => n8328);
   U5140 : OAI22_X1 port map( A1 => n20434, A2 => n19969, B1 => n4216, B2 => 
                           n19980, ZN => n8329);
   U5141 : OAI22_X1 port map( A1 => n20437, A2 => n19969, B1 => n4215, B2 => 
                           n19980, ZN => n8330);
   U5142 : OAI22_X1 port map( A1 => n20440, A2 => n19968, B1 => n4214, B2 => 
                           n19979, ZN => n8331);
   U5143 : OAI22_X1 port map( A1 => n20443, A2 => n19968, B1 => n4213, B2 => 
                           n19979, ZN => n8332);
   U5144 : OAI22_X1 port map( A1 => n20446, A2 => n19968, B1 => n4212, B2 => 
                           n19979, ZN => n8333);
   U5145 : OAI22_X1 port map( A1 => n20449, A2 => n19968, B1 => n4211, B2 => 
                           n19979, ZN => n8334);
   U5146 : OAI22_X1 port map( A1 => n20452, A2 => n19968, B1 => n4210, B2 => 
                           n19978, ZN => n8335);
   U5147 : OAI22_X1 port map( A1 => n20455, A2 => n19968, B1 => n4209, B2 => 
                           n19978, ZN => n8336);
   U5148 : OAI22_X1 port map( A1 => n20458, A2 => n19968, B1 => n4208, B2 => 
                           n19978, ZN => n8337);
   U5149 : OAI22_X1 port map( A1 => n20461, A2 => n19968, B1 => n4207, B2 => 
                           n19978, ZN => n8338);
   U5150 : OAI22_X1 port map( A1 => n20464, A2 => n19968, B1 => n4206, B2 => 
                           n19977, ZN => n8339);
   U5151 : OAI22_X1 port map( A1 => n20467, A2 => n19968, B1 => n4205, B2 => 
                           n19977, ZN => n8340);
   U5152 : OAI22_X1 port map( A1 => n20470, A2 => n19968, B1 => n4204, B2 => 
                           n19977, ZN => n8341);
   U5153 : OAI22_X1 port map( A1 => n20473, A2 => n19968, B1 => n4203, B2 => 
                           n19977, ZN => n8342);
   U5154 : OAI22_X1 port map( A1 => n20476, A2 => n19970, B1 => n4202, B2 => 
                           n19976, ZN => n8343);
   U5155 : OAI22_X1 port map( A1 => n20479, A2 => n19969, B1 => n4201, B2 => 
                           n19976, ZN => n8344);
   U5156 : OAI22_X1 port map( A1 => n20482, A2 => n19968, B1 => n4200, B2 => 
                           n19976, ZN => n8345);
   U5157 : OAI22_X1 port map( A1 => n20485, A2 => n19970, B1 => n4199, B2 => 
                           n19976, ZN => n8346);
   U5158 : OAI22_X1 port map( A1 => n20488, A2 => n19969, B1 => n4198, B2 => 
                           n19975, ZN => n8347);
   U5159 : OAI22_X1 port map( A1 => n20491, A2 => n19968, B1 => n4197, B2 => 
                           n19975, ZN => n8348);
   U5160 : OAI22_X1 port map( A1 => n20494, A2 => n19970, B1 => n4196, B2 => 
                           n19975, ZN => n8349);
   U5161 : OAI22_X1 port map( A1 => n20497, A2 => n19969, B1 => n4195, B2 => 
                           n19975, ZN => n8350);
   U5162 : OAI22_X1 port map( A1 => n20500, A2 => n19968, B1 => n4194, B2 => 
                           n19974, ZN => n8351);
   U5163 : OAI22_X1 port map( A1 => n20503, A2 => n19970, B1 => n4193, B2 => 
                           n19974, ZN => n8352);
   U5164 : OAI22_X1 port map( A1 => n20506, A2 => n19969, B1 => n4192, B2 => 
                           n19974, ZN => n8353);
   U5165 : OAI22_X1 port map( A1 => n20509, A2 => n19969, B1 => n4191, B2 => 
                           n19974, ZN => n8354);
   U5166 : OAI22_X1 port map( A1 => n20512, A2 => n19970, B1 => n4190, B2 => 
                           n19973, ZN => n8355);
   U5167 : OAI22_X1 port map( A1 => n20515, A2 => n19969, B1 => n4189, B2 => 
                           n19973, ZN => n8356);
   U5168 : OAI22_X1 port map( A1 => n20518, A2 => n19968, B1 => n4188, B2 => 
                           n19973, ZN => n8357);
   U5169 : OAI22_X1 port map( A1 => n20521, A2 => n19968, B1 => n4187, B2 => 
                           n19973, ZN => n8358);
   U5170 : OAI22_X1 port map( A1 => n20524, A2 => n19970, B1 => n4186, B2 => 
                           n19972, ZN => n8359);
   U5171 : OAI22_X1 port map( A1 => n20527, A2 => n19969, B1 => n4185, B2 => 
                           n19972, ZN => n8360);
   U5172 : OAI22_X1 port map( A1 => n20530, A2 => n19968, B1 => n4184, B2 => 
                           n19972, ZN => n8361);
   U5173 : OAI22_X1 port map( A1 => n20533, A2 => n19970, B1 => n4183, B2 => 
                           n19972, ZN => n8362);
   U5174 : OAI22_X1 port map( A1 => n20536, A2 => n19970, B1 => n4182, B2 => 
                           n19971, ZN => n8363);
   U5175 : OAI22_X1 port map( A1 => n20539, A2 => n19969, B1 => n4181, B2 => 
                           n19971, ZN => n8364);
   U5176 : OAI22_X1 port map( A1 => n20542, A2 => n19968, B1 => n4180, B2 => 
                           n19971, ZN => n8365);
   U5177 : OAI22_X1 port map( A1 => n20573, A2 => n19969, B1 => n4179, B2 => 
                           n19971, ZN => n8366);
   U5178 : OAI22_X1 port map( A1 => n20356, A2 => n19969, B1 => n4242, B2 => 
                           n19986, ZN => n8303);
   U5179 : OAI22_X1 port map( A1 => n20359, A2 => n19968, B1 => n4241, B2 => 
                           n19986, ZN => n8304);
   U5180 : OAI22_X1 port map( A1 => n20362, A2 => n19968, B1 => n4240, B2 => 
                           n19986, ZN => n8305);
   U5181 : OAI22_X1 port map( A1 => n20365, A2 => n19970, B1 => n4239, B2 => 
                           n19986, ZN => n8306);
   U5182 : OAI22_X1 port map( A1 => n20368, A2 => n19830, B1 => n4576, B2 => 
                           n19845, ZN => n7987);
   U5183 : OAI22_X1 port map( A1 => n20371, A2 => n19830, B1 => n4575, B2 => 
                           n19845, ZN => n7988);
   U5184 : OAI22_X1 port map( A1 => n20374, A2 => n19830, B1 => n4574, B2 => 
                           n19845, ZN => n7989);
   U5185 : OAI22_X1 port map( A1 => n20377, A2 => n19830, B1 => n4573, B2 => 
                           n19845, ZN => n7990);
   U5186 : OAI22_X1 port map( A1 => n20380, A2 => n19830, B1 => n4572, B2 => 
                           n19844, ZN => n7991);
   U5187 : OAI22_X1 port map( A1 => n20383, A2 => n19830, B1 => n4571, B2 => 
                           n19844, ZN => n7992);
   U5188 : OAI22_X1 port map( A1 => n20386, A2 => n19830, B1 => n4570, B2 => 
                           n19844, ZN => n7993);
   U5189 : OAI22_X1 port map( A1 => n20389, A2 => n19830, B1 => n4569, B2 => 
                           n19844, ZN => n7994);
   U5190 : OAI22_X1 port map( A1 => n20392, A2 => n19830, B1 => n4568, B2 => 
                           n19843, ZN => n7995);
   U5191 : OAI22_X1 port map( A1 => n20395, A2 => n19830, B1 => n4567, B2 => 
                           n19843, ZN => n7996);
   U5192 : OAI22_X1 port map( A1 => n20398, A2 => n19830, B1 => n4566, B2 => 
                           n19843, ZN => n7997);
   U5193 : OAI22_X1 port map( A1 => n20401, A2 => n19830, B1 => n4565, B2 => 
                           n19843, ZN => n7998);
   U5194 : OAI22_X1 port map( A1 => n20404, A2 => n19829, B1 => n4564, B2 => 
                           n19842, ZN => n7999);
   U5195 : OAI22_X1 port map( A1 => n20407, A2 => n19829, B1 => n4563, B2 => 
                           n19842, ZN => n8000);
   U5196 : OAI22_X1 port map( A1 => n20410, A2 => n19829, B1 => n4562, B2 => 
                           n19842, ZN => n8001);
   U5197 : OAI22_X1 port map( A1 => n20413, A2 => n19829, B1 => n4561, B2 => 
                           n19842, ZN => n8002);
   U5198 : OAI22_X1 port map( A1 => n20416, A2 => n19829, B1 => n4560, B2 => 
                           n19841, ZN => n8003);
   U5199 : OAI22_X1 port map( A1 => n20419, A2 => n19829, B1 => n4559, B2 => 
                           n19841, ZN => n8004);
   U5200 : OAI22_X1 port map( A1 => n20422, A2 => n19829, B1 => n4558, B2 => 
                           n19841, ZN => n8005);
   U5201 : OAI22_X1 port map( A1 => n20425, A2 => n19829, B1 => n4557, B2 => 
                           n19841, ZN => n8006);
   U5202 : OAI22_X1 port map( A1 => n20428, A2 => n19829, B1 => n4556, B2 => 
                           n19840, ZN => n8007);
   U5203 : OAI22_X1 port map( A1 => n20431, A2 => n19829, B1 => n4555, B2 => 
                           n19840, ZN => n8008);
   U5204 : OAI22_X1 port map( A1 => n20434, A2 => n19829, B1 => n4554, B2 => 
                           n19840, ZN => n8009);
   U5205 : OAI22_X1 port map( A1 => n20437, A2 => n19829, B1 => n4553, B2 => 
                           n19840, ZN => n8010);
   U5206 : OAI22_X1 port map( A1 => n20440, A2 => n19828, B1 => n4552, B2 => 
                           n19839, ZN => n8011);
   U5207 : OAI22_X1 port map( A1 => n20443, A2 => n19828, B1 => n4551, B2 => 
                           n19839, ZN => n8012);
   U5208 : OAI22_X1 port map( A1 => n20446, A2 => n19828, B1 => n4550, B2 => 
                           n19839, ZN => n8013);
   U5209 : OAI22_X1 port map( A1 => n20449, A2 => n19828, B1 => n4549, B2 => 
                           n19839, ZN => n8014);
   U5210 : OAI22_X1 port map( A1 => n20452, A2 => n19828, B1 => n4548, B2 => 
                           n19838, ZN => n8015);
   U5211 : OAI22_X1 port map( A1 => n20455, A2 => n19828, B1 => n4547, B2 => 
                           n19838, ZN => n8016);
   U5212 : OAI22_X1 port map( A1 => n20458, A2 => n19828, B1 => n4546, B2 => 
                           n19838, ZN => n8017);
   U5213 : OAI22_X1 port map( A1 => n20461, A2 => n19828, B1 => n4545, B2 => 
                           n19838, ZN => n8018);
   U5214 : OAI22_X1 port map( A1 => n20464, A2 => n19828, B1 => n4544, B2 => 
                           n19837, ZN => n8019);
   U5215 : OAI22_X1 port map( A1 => n20467, A2 => n19828, B1 => n4543, B2 => 
                           n19837, ZN => n8020);
   U5216 : OAI22_X1 port map( A1 => n20470, A2 => n19828, B1 => n4542, B2 => 
                           n19837, ZN => n8021);
   U5217 : OAI22_X1 port map( A1 => n20473, A2 => n19828, B1 => n4541, B2 => 
                           n19837, ZN => n8022);
   U5218 : OAI22_X1 port map( A1 => n20476, A2 => n19830, B1 => n4540, B2 => 
                           n19836, ZN => n8023);
   U5219 : OAI22_X1 port map( A1 => n20479, A2 => n19829, B1 => n4539, B2 => 
                           n19836, ZN => n8024);
   U5220 : OAI22_X1 port map( A1 => n20482, A2 => n19828, B1 => n4538, B2 => 
                           n19836, ZN => n8025);
   U5221 : OAI22_X1 port map( A1 => n20485, A2 => n19830, B1 => n4537, B2 => 
                           n19836, ZN => n8026);
   U5222 : OAI22_X1 port map( A1 => n20488, A2 => n19829, B1 => n4536, B2 => 
                           n19835, ZN => n8027);
   U5223 : OAI22_X1 port map( A1 => n20491, A2 => n19828, B1 => n4535, B2 => 
                           n19835, ZN => n8028);
   U5224 : OAI22_X1 port map( A1 => n20494, A2 => n19830, B1 => n4534, B2 => 
                           n19835, ZN => n8029);
   U5225 : OAI22_X1 port map( A1 => n20497, A2 => n19829, B1 => n4533, B2 => 
                           n19835, ZN => n8030);
   U5226 : OAI22_X1 port map( A1 => n20500, A2 => n19828, B1 => n4532, B2 => 
                           n19834, ZN => n8031);
   U5227 : OAI22_X1 port map( A1 => n20503, A2 => n19830, B1 => n4531, B2 => 
                           n19834, ZN => n8032);
   U5228 : OAI22_X1 port map( A1 => n20506, A2 => n19829, B1 => n4530, B2 => 
                           n19834, ZN => n8033);
   U5229 : OAI22_X1 port map( A1 => n20509, A2 => n19829, B1 => n4529, B2 => 
                           n19834, ZN => n8034);
   U5230 : OAI22_X1 port map( A1 => n20512, A2 => n19830, B1 => n4528, B2 => 
                           n19833, ZN => n8035);
   U5231 : OAI22_X1 port map( A1 => n20515, A2 => n19829, B1 => n4527, B2 => 
                           n19833, ZN => n8036);
   U5232 : OAI22_X1 port map( A1 => n20518, A2 => n19828, B1 => n4526, B2 => 
                           n19833, ZN => n8037);
   U5233 : OAI22_X1 port map( A1 => n20521, A2 => n19828, B1 => n4525, B2 => 
                           n19833, ZN => n8038);
   U5234 : OAI22_X1 port map( A1 => n20524, A2 => n19830, B1 => n4524, B2 => 
                           n19832, ZN => n8039);
   U5235 : OAI22_X1 port map( A1 => n20527, A2 => n19829, B1 => n4523, B2 => 
                           n19832, ZN => n8040);
   U5236 : OAI22_X1 port map( A1 => n20530, A2 => n19828, B1 => n4522, B2 => 
                           n19832, ZN => n8041);
   U5237 : OAI22_X1 port map( A1 => n20533, A2 => n19830, B1 => n4521, B2 => 
                           n19832, ZN => n8042);
   U5238 : OAI22_X1 port map( A1 => n20536, A2 => n19830, B1 => n4520, B2 => 
                           n19831, ZN => n8043);
   U5239 : OAI22_X1 port map( A1 => n20539, A2 => n19829, B1 => n4519, B2 => 
                           n19831, ZN => n8044);
   U5240 : OAI22_X1 port map( A1 => n20542, A2 => n19828, B1 => n4518, B2 => 
                           n19831, ZN => n8045);
   U5241 : OAI22_X1 port map( A1 => n20573, A2 => n19829, B1 => n4517, B2 => 
                           n19831, ZN => n8046);
   U5242 : OAI22_X1 port map( A1 => n20356, A2 => n19829, B1 => n4580, B2 => 
                           n19846, ZN => n7983);
   U5243 : OAI22_X1 port map( A1 => n20359, A2 => n19828, B1 => n4579, B2 => 
                           n19846, ZN => n7984);
   U5244 : OAI22_X1 port map( A1 => n20362, A2 => n19828, B1 => n4578, B2 => 
                           n19846, ZN => n7985);
   U5245 : OAI22_X1 port map( A1 => n20365, A2 => n19830, B1 => n4577, B2 => 
                           n19846, ZN => n7986);
   U5246 : AOI22_X1 port map( A1 => n18993, A2 => n6751, B1 => n18987, B2 => 
                           registers_14_39_port, ZN => n6750);
   U5247 : AOI22_X1 port map( A1 => n18993, A2 => n6683, B1 => n18987, B2 => 
                           registers_14_40_port, ZN => n6682);
   U5248 : AOI22_X1 port map( A1 => n18993, A2 => n6616, B1 => n18987, B2 => 
                           registers_14_41_port, ZN => n6615);
   U5249 : AOI22_X1 port map( A1 => n18993, A2 => n6550, B1 => n18987, B2 => 
                           registers_14_42_port, ZN => n6549);
   U5250 : AOI22_X1 port map( A1 => n18993, A2 => n6484, B1 => n18987, B2 => 
                           registers_14_43_port, ZN => n6483);
   U5251 : AOI22_X1 port map( A1 => n18993, A2 => n6418, B1 => n18987, B2 => 
                           registers_14_44_port, ZN => n6417);
   U5252 : AOI22_X1 port map( A1 => n18993, A2 => n6352, B1 => n18987, B2 => 
                           registers_14_45_port, ZN => n6351);
   U5253 : AOI22_X1 port map( A1 => n18993, A2 => n6286, B1 => n18987, B2 => 
                           registers_14_46_port, ZN => n6285);
   U5254 : AOI22_X1 port map( A1 => n18993, A2 => n6220, B1 => n18987, B2 => 
                           registers_14_47_port, ZN => n6219);
   U5255 : AOI22_X1 port map( A1 => n18994, A2 => n6154, B1 => n18988, B2 => 
                           registers_14_48_port, ZN => n6153);
   U5256 : AOI22_X1 port map( A1 => n18994, A2 => n6088, B1 => n18988, B2 => 
                           registers_14_49_port, ZN => n6087);
   U5257 : AOI22_X1 port map( A1 => n18994, A2 => n6020, B1 => n18988, B2 => 
                           registers_14_50_port, ZN => n6019);
   U5258 : AOI22_X1 port map( A1 => n18994, A2 => n5952, B1 => n18988, B2 => 
                           registers_14_51_port, ZN => n5951);
   U5259 : AOI22_X1 port map( A1 => n18994, A2 => n5885, B1 => n18988, B2 => 
                           registers_14_52_port, ZN => n5884);
   U5260 : AOI22_X1 port map( A1 => n18994, A2 => n5818, B1 => n18988, B2 => 
                           registers_14_53_port, ZN => n5817);
   U5261 : AOI22_X1 port map( A1 => n18994, A2 => n5746, B1 => n18988, B2 => 
                           registers_14_54_port, ZN => n5745);
   U5262 : AOI22_X1 port map( A1 => n18994, A2 => n5676, B1 => n18988, B2 => 
                           registers_14_55_port, ZN => n5675);
   U5263 : AOI22_X1 port map( A1 => n18994, A2 => n5608, B1 => n18988, B2 => 
                           registers_14_56_port, ZN => n5607);
   U5264 : AOI22_X1 port map( A1 => n18994, A2 => n5539, B1 => n18988, B2 => 
                           registers_14_57_port, ZN => n5538);
   U5265 : AOI22_X1 port map( A1 => n18994, A2 => n5470, B1 => n18988, B2 => 
                           registers_14_58_port, ZN => n5469);
   U5266 : AOI22_X1 port map( A1 => n18994, A2 => n5402, B1 => n18988, B2 => 
                           registers_14_59_port, ZN => n5401);
   U5267 : AOI22_X1 port map( A1 => n18990, A2 => n11690, B1 => n18984, B2 => 
                           registers_14_0_port, ZN => n11689);
   U5268 : AOI22_X1 port map( A1 => n18990, A2 => n11546, B1 => n18984, B2 => 
                           registers_14_1_port, ZN => n11545);
   U5269 : AOI22_X1 port map( A1 => n18990, A2 => n11478, B1 => n18984, B2 => 
                           registers_14_2_port, ZN => n11477);
   U5270 : AOI22_X1 port map( A1 => n18990, A2 => n11411, B1 => n18984, B2 => 
                           registers_14_3_port, ZN => n11410);
   U5271 : AOI22_X1 port map( A1 => n18990, A2 => n11344, B1 => n18984, B2 => 
                           registers_14_4_port, ZN => n11343);
   U5272 : AOI22_X1 port map( A1 => n18990, A2 => n11276, B1 => n18984, B2 => 
                           registers_14_5_port, ZN => n11275);
   U5273 : AOI22_X1 port map( A1 => n18990, A2 => n11209, B1 => n18984, B2 => 
                           registers_14_6_port, ZN => n11208);
   U5274 : AOI22_X1 port map( A1 => n18990, A2 => n11142, B1 => n18984, B2 => 
                           registers_14_7_port, ZN => n11141);
   U5275 : AOI22_X1 port map( A1 => n18990, A2 => n11075, B1 => n18984, B2 => 
                           registers_14_8_port, ZN => n11074);
   U5276 : AOI22_X1 port map( A1 => n18990, A2 => n11007, B1 => n18984, B2 => 
                           registers_14_9_port, ZN => n11006);
   U5277 : AOI22_X1 port map( A1 => n18990, A2 => n10940, B1 => n18984, B2 => 
                           registers_14_10_port, ZN => n10939);
   U5278 : AOI22_X1 port map( A1 => n18990, A2 => n10873, B1 => n18984, B2 => 
                           registers_14_11_port, ZN => n10872);
   U5279 : AOI22_X1 port map( A1 => n18991, A2 => n10806, B1 => n18985, B2 => 
                           registers_14_12_port, ZN => n10805);
   U5280 : AOI22_X1 port map( A1 => n18991, A2 => n10738, B1 => n18985, B2 => 
                           registers_14_13_port, ZN => n10737);
   U5281 : AOI22_X1 port map( A1 => n18991, A2 => n10671, B1 => n18985, B2 => 
                           registers_14_14_port, ZN => n10670);
   U5282 : AOI22_X1 port map( A1 => n18991, A2 => n10604, B1 => n18985, B2 => 
                           registers_14_15_port, ZN => n10603);
   U5283 : AOI22_X1 port map( A1 => n18991, A2 => n10537, B1 => n18985, B2 => 
                           registers_14_16_port, ZN => n10535);
   U5284 : AOI22_X1 port map( A1 => n18991, A2 => n10469, B1 => n18985, B2 => 
                           registers_14_17_port, ZN => n10468);
   U5285 : AOI22_X1 port map( A1 => n18991, A2 => n10402, B1 => n18985, B2 => 
                           registers_14_18_port, ZN => n10401);
   U5286 : AOI22_X1 port map( A1 => n18991, A2 => n10335, B1 => n18985, B2 => 
                           registers_14_19_port, ZN => n10334);
   U5287 : AOI22_X1 port map( A1 => n18991, A2 => n10267, B1 => n18985, B2 => 
                           registers_14_20_port, ZN => n10266);
   U5288 : AOI22_X1 port map( A1 => n18991, A2 => n10200, B1 => n18985, B2 => 
                           registers_14_21_port, ZN => n10199);
   U5289 : AOI22_X1 port map( A1 => n18991, A2 => n10133, B1 => n18985, B2 => 
                           registers_14_22_port, ZN => n10132);
   U5290 : AOI22_X1 port map( A1 => n18991, A2 => n10066, B1 => n18985, B2 => 
                           registers_14_23_port, ZN => n10065);
   U5291 : AOI22_X1 port map( A1 => n18992, A2 => n9998, B1 => n18986, B2 => 
                           registers_14_24_port, ZN => n9997);
   U5292 : AOI22_X1 port map( A1 => n18992, A2 => n9931, B1 => n18986, B2 => 
                           registers_14_25_port, ZN => n9930);
   U5293 : AOI22_X1 port map( A1 => n18992, A2 => n9864, B1 => n18986, B2 => 
                           registers_14_26_port, ZN => n9863);
   U5294 : AOI22_X1 port map( A1 => n18992, A2 => n9797, B1 => n18986, B2 => 
                           registers_14_27_port, ZN => n9796);
   U5295 : AOI22_X1 port map( A1 => n18992, A2 => n9729, B1 => n18986, B2 => 
                           registers_14_28_port, ZN => n9728);
   U5296 : AOI22_X1 port map( A1 => n18992, A2 => n9662, B1 => n18986, B2 => 
                           registers_14_29_port, ZN => n9661);
   U5297 : AOI22_X1 port map( A1 => n18992, A2 => n9595, B1 => n18986, B2 => 
                           registers_14_30_port, ZN => n9594);
   U5298 : AOI22_X1 port map( A1 => n18992, A2 => n9527, B1 => n18986, B2 => 
                           registers_14_31_port, ZN => n9526);
   U5299 : AOI22_X1 port map( A1 => n18992, A2 => n9460, B1 => n18986, B2 => 
                           registers_14_32_port, ZN => n9459);
   U5300 : AOI22_X1 port map( A1 => n18992, A2 => n9393, B1 => n18986, B2 => 
                           registers_14_33_port, ZN => n9392);
   U5301 : AOI22_X1 port map( A1 => n18992, A2 => n9326, B1 => n18986, B2 => 
                           registers_14_34_port, ZN => n9325);
   U5302 : AOI22_X1 port map( A1 => n18992, A2 => n7018, B1 => n18986, B2 => 
                           registers_14_35_port, ZN => n7017);
   U5303 : AOI22_X1 port map( A1 => n18995, A2 => n5332, B1 => n18989, B2 => 
                           registers_14_60_port, ZN => n5331);
   U5304 : AOI22_X1 port map( A1 => n18995, A2 => n4719, B1 => n18989, B2 => 
                           registers_14_61_port, ZN => n4718);
   U5305 : AOI22_X1 port map( A1 => n18995, A2 => n3437, B1 => n18989, B2 => 
                           registers_14_62_port, ZN => n3436);
   U5306 : AOI22_X1 port map( A1 => n18995, A2 => n3164, B1 => n18989, B2 => 
                           registers_14_63_port, ZN => n3162);
   U5307 : AOI22_X1 port map( A1 => n18993, A2 => n6952, B1 => n18987, B2 => 
                           registers_14_36_port, ZN => n6951);
   U5308 : AOI22_X1 port map( A1 => n18993, A2 => n6885, B1 => n18987, B2 => 
                           registers_14_37_port, ZN => n6884);
   U5309 : OAI22_X1 port map( A1 => n20367, A2 => n19522, B1 => n5835, B2 => 
                           n19537, ZN => n7283);
   U5310 : OAI22_X1 port map( A1 => n20370, A2 => n19522, B1 => n5769, B2 => 
                           n19537, ZN => n7284);
   U5311 : OAI22_X1 port map( A1 => n20373, A2 => n19522, B1 => n5767, B2 => 
                           n19537, ZN => n7285);
   U5312 : OAI22_X1 port map( A1 => n20376, A2 => n19522, B1 => n5766, B2 => 
                           n19537, ZN => n7286);
   U5313 : OAI22_X1 port map( A1 => n20379, A2 => n19522, B1 => n5765, B2 => 
                           n19536, ZN => n7287);
   U5314 : OAI22_X1 port map( A1 => n20382, A2 => n19522, B1 => n5764, B2 => 
                           n19536, ZN => n7288);
   U5315 : OAI22_X1 port map( A1 => n20385, A2 => n19522, B1 => n5763, B2 => 
                           n19536, ZN => n7289);
   U5316 : OAI22_X1 port map( A1 => n20388, A2 => n19522, B1 => n5698, B2 => 
                           n19536, ZN => n7290);
   U5317 : OAI22_X1 port map( A1 => n20391, A2 => n19522, B1 => n5696, B2 => 
                           n19535, ZN => n7291);
   U5318 : OAI22_X1 port map( A1 => n20394, A2 => n19522, B1 => n5695, B2 => 
                           n19535, ZN => n7292);
   U5319 : OAI22_X1 port map( A1 => n20397, A2 => n19522, B1 => n5694, B2 => 
                           n19535, ZN => n7293);
   U5320 : OAI22_X1 port map( A1 => n20400, A2 => n19522, B1 => n5629, B2 => 
                           n19535, ZN => n7294);
   U5321 : OAI22_X1 port map( A1 => n20403, A2 => n19521, B1 => n5627, B2 => 
                           n19534, ZN => n7295);
   U5322 : OAI22_X1 port map( A1 => n20406, A2 => n19521, B1 => n5562, B2 => 
                           n19534, ZN => n7296);
   U5323 : OAI22_X1 port map( A1 => n20409, A2 => n19521, B1 => n5560, B2 => 
                           n19534, ZN => n7297);
   U5324 : OAI22_X1 port map( A1 => n20412, A2 => n19521, B1 => n5559, B2 => 
                           n19534, ZN => n7298);
   U5325 : OAI22_X1 port map( A1 => n20415, A2 => n19521, B1 => n5494, B2 => 
                           n19533, ZN => n7299);
   U5326 : OAI22_X1 port map( A1 => n20418, A2 => n19521, B1 => n5492, B2 => 
                           n19533, ZN => n7300);
   U5327 : OAI22_X1 port map( A1 => n20421, A2 => n19521, B1 => n5491, B2 => 
                           n19533, ZN => n7301);
   U5328 : OAI22_X1 port map( A1 => n20424, A2 => n19521, B1 => n5426, B2 => 
                           n19533, ZN => n7302);
   U5329 : OAI22_X1 port map( A1 => n20427, A2 => n19521, B1 => n5424, B2 => 
                           n19532, ZN => n7303);
   U5330 : OAI22_X1 port map( A1 => n20430, A2 => n19521, B1 => n5359, B2 => 
                           n19532, ZN => n7304);
   U5331 : OAI22_X1 port map( A1 => n20433, A2 => n19521, B1 => n5357, B2 => 
                           n19532, ZN => n7305);
   U5332 : OAI22_X1 port map( A1 => n20436, A2 => n19521, B1 => n5356, B2 => 
                           n19532, ZN => n7306);
   U5333 : OAI22_X1 port map( A1 => n20439, A2 => n19522, B1 => n5355, B2 => 
                           n19531, ZN => n7307);
   U5334 : OAI22_X1 port map( A1 => n20442, A2 => n19521, B1 => n5291, B2 => 
                           n19531, ZN => n7308);
   U5335 : OAI22_X1 port map( A1 => n20445, A2 => n19520, B1 => n5290, B2 => 
                           n19531, ZN => n7309);
   U5336 : OAI22_X1 port map( A1 => n20448, A2 => n19522, B1 => n5289, B2 => 
                           n19531, ZN => n7310);
   U5337 : OAI22_X1 port map( A1 => n20451, A2 => n19521, B1 => n5288, B2 => 
                           n19530, ZN => n7311);
   U5338 : OAI22_X1 port map( A1 => n20454, A2 => n19520, B1 => n5287, B2 => 
                           n19530, ZN => n7312);
   U5339 : OAI22_X1 port map( A1 => n20457, A2 => n19522, B1 => n5286, B2 => 
                           n19530, ZN => n7313);
   U5340 : OAI22_X1 port map( A1 => n20460, A2 => n19521, B1 => n5285, B2 => 
                           n19530, ZN => n7314);
   U5341 : OAI22_X1 port map( A1 => n20463, A2 => n19520, B1 => n5284, B2 => 
                           n19529, ZN => n7315);
   U5342 : OAI22_X1 port map( A1 => n20466, A2 => n19522, B1 => n5283, B2 => 
                           n19529, ZN => n7316);
   U5343 : OAI22_X1 port map( A1 => n20472, A2 => n19521, B1 => n5281, B2 => 
                           n19529, ZN => n7318);
   U5344 : OAI22_X1 port map( A1 => n20475, A2 => n19520, B1 => n5280, B2 => 
                           n19528, ZN => n7319);
   U5345 : OAI22_X1 port map( A1 => n20478, A2 => n19520, B1 => n5279, B2 => 
                           n19528, ZN => n7320);
   U5346 : OAI22_X1 port map( A1 => n20481, A2 => n19520, B1 => n5278, B2 => 
                           n19528, ZN => n7321);
   U5347 : OAI22_X1 port map( A1 => n20484, A2 => n19520, B1 => n5277, B2 => 
                           n19528, ZN => n7322);
   U5348 : OAI22_X1 port map( A1 => n20487, A2 => n19520, B1 => n5276, B2 => 
                           n19527, ZN => n7323);
   U5349 : OAI22_X1 port map( A1 => n20490, A2 => n19520, B1 => n5275, B2 => 
                           n19527, ZN => n7324);
   U5350 : OAI22_X1 port map( A1 => n20493, A2 => n19520, B1 => n5274, B2 => 
                           n19527, ZN => n7325);
   U5351 : OAI22_X1 port map( A1 => n20496, A2 => n19520, B1 => n5273, B2 => 
                           n19527, ZN => n7326);
   U5352 : OAI22_X1 port map( A1 => n20499, A2 => n19520, B1 => n5272, B2 => 
                           n19526, ZN => n7327);
   U5353 : OAI22_X1 port map( A1 => n20502, A2 => n19520, B1 => n5271, B2 => 
                           n19526, ZN => n7328);
   U5354 : OAI22_X1 port map( A1 => n20505, A2 => n19520, B1 => n5270, B2 => 
                           n19526, ZN => n7329);
   U5355 : OAI22_X1 port map( A1 => n20508, A2 => n19520, B1 => n5269, B2 => 
                           n19526, ZN => n7330);
   U5356 : OAI22_X1 port map( A1 => n20511, A2 => n19522, B1 => n5268, B2 => 
                           n19525, ZN => n7331);
   U5357 : OAI22_X1 port map( A1 => n20514, A2 => n19521, B1 => n5267, B2 => 
                           n19525, ZN => n7332);
   U5358 : OAI22_X1 port map( A1 => n20517, A2 => n19520, B1 => n5266, B2 => 
                           n19525, ZN => n7333);
   U5359 : OAI22_X1 port map( A1 => n20520, A2 => n19520, B1 => n5265, B2 => 
                           n19525, ZN => n7334);
   U5360 : OAI22_X1 port map( A1 => n20523, A2 => n19522, B1 => n5264, B2 => 
                           n19524, ZN => n7335);
   U5361 : OAI22_X1 port map( A1 => n20526, A2 => n19521, B1 => n5263, B2 => 
                           n19524, ZN => n7336);
   U5362 : OAI22_X1 port map( A1 => n20529, A2 => n19522, B1 => n5262, B2 => 
                           n19524, ZN => n7337);
   U5363 : OAI22_X1 port map( A1 => n20532, A2 => n19520, B1 => n5261, B2 => 
                           n19524, ZN => n7338);
   U5364 : OAI22_X1 port map( A1 => n20535, A2 => n19522, B1 => n5260, B2 => 
                           n19523, ZN => n7339);
   U5365 : OAI22_X1 port map( A1 => n20538, A2 => n19521, B1 => n5259, B2 => 
                           n19523, ZN => n7340);
   U5366 : OAI22_X1 port map( A1 => n20541, A2 => n19521, B1 => n5258, B2 => 
                           n19523, ZN => n7341);
   U5367 : OAI22_X1 port map( A1 => n20572, A2 => n19520, B1 => n5257, B2 => 
                           n19523, ZN => n7342);
   U5368 : OAI22_X1 port map( A1 => n20355, A2 => n19521, B1 => n6033, B2 => 
                           n19538, ZN => n7279);
   U5369 : OAI22_X1 port map( A1 => n20358, A2 => n19520, B1 => n5968, B2 => 
                           n19538, ZN => n7280);
   U5370 : OAI22_X1 port map( A1 => n20361, A2 => n19520, B1 => n5966, B2 => 
                           n19538, ZN => n7281);
   U5371 : OAI22_X1 port map( A1 => n20364, A2 => n19522, B1 => n5901, B2 => 
                           n19538, ZN => n7282);
   U5372 : OAI22_X1 port map( A1 => n20367, A2 => n19718, B1 => n4846, B2 => 
                           n19733, ZN => n7731);
   U5373 : OAI22_X1 port map( A1 => n20370, A2 => n19718, B1 => n4845, B2 => 
                           n19733, ZN => n7732);
   U5374 : OAI22_X1 port map( A1 => n20373, A2 => n19718, B1 => n4844, B2 => 
                           n19733, ZN => n7733);
   U5375 : OAI22_X1 port map( A1 => n20376, A2 => n19718, B1 => n4843, B2 => 
                           n19733, ZN => n7734);
   U5376 : OAI22_X1 port map( A1 => n20379, A2 => n19718, B1 => n4842, B2 => 
                           n19732, ZN => n7735);
   U5377 : OAI22_X1 port map( A1 => n20382, A2 => n19718, B1 => n4841, B2 => 
                           n19732, ZN => n7736);
   U5378 : OAI22_X1 port map( A1 => n20385, A2 => n19718, B1 => n4840, B2 => 
                           n19732, ZN => n7737);
   U5379 : OAI22_X1 port map( A1 => n20388, A2 => n19718, B1 => n4839, B2 => 
                           n19732, ZN => n7738);
   U5380 : OAI22_X1 port map( A1 => n20391, A2 => n19718, B1 => n4838, B2 => 
                           n19731, ZN => n7739);
   U5381 : OAI22_X1 port map( A1 => n20394, A2 => n19718, B1 => n4837, B2 => 
                           n19731, ZN => n7740);
   U5382 : OAI22_X1 port map( A1 => n20397, A2 => n19718, B1 => n4836, B2 => 
                           n19731, ZN => n7741);
   U5383 : OAI22_X1 port map( A1 => n20400, A2 => n19718, B1 => n4835, B2 => 
                           n19731, ZN => n7742);
   U5384 : OAI22_X1 port map( A1 => n20403, A2 => n19717, B1 => n4834, B2 => 
                           n19730, ZN => n7743);
   U5385 : OAI22_X1 port map( A1 => n20406, A2 => n19717, B1 => n4833, B2 => 
                           n19730, ZN => n7744);
   U5386 : OAI22_X1 port map( A1 => n20409, A2 => n19717, B1 => n4832, B2 => 
                           n19730, ZN => n7745);
   U5387 : OAI22_X1 port map( A1 => n20412, A2 => n19717, B1 => n4831, B2 => 
                           n19730, ZN => n7746);
   U5388 : OAI22_X1 port map( A1 => n20415, A2 => n19717, B1 => n4830, B2 => 
                           n19729, ZN => n7747);
   U5389 : OAI22_X1 port map( A1 => n20418, A2 => n19717, B1 => n4829, B2 => 
                           n19729, ZN => n7748);
   U5390 : OAI22_X1 port map( A1 => n20421, A2 => n19717, B1 => n4828, B2 => 
                           n19729, ZN => n7749);
   U5391 : OAI22_X1 port map( A1 => n20424, A2 => n19717, B1 => n4827, B2 => 
                           n19729, ZN => n7750);
   U5392 : OAI22_X1 port map( A1 => n20427, A2 => n19717, B1 => n4826, B2 => 
                           n19728, ZN => n7751);
   U5393 : OAI22_X1 port map( A1 => n20430, A2 => n19717, B1 => n4825, B2 => 
                           n19728, ZN => n7752);
   U5394 : OAI22_X1 port map( A1 => n20433, A2 => n19717, B1 => n4824, B2 => 
                           n19728, ZN => n7753);
   U5395 : OAI22_X1 port map( A1 => n20436, A2 => n19717, B1 => n4823, B2 => 
                           n19728, ZN => n7754);
   U5396 : OAI22_X1 port map( A1 => n20439, A2 => n19716, B1 => n4822, B2 => 
                           n19727, ZN => n7755);
   U5397 : OAI22_X1 port map( A1 => n20442, A2 => n19716, B1 => n4821, B2 => 
                           n19727, ZN => n7756);
   U5398 : OAI22_X1 port map( A1 => n20445, A2 => n19716, B1 => n4820, B2 => 
                           n19727, ZN => n7757);
   U5399 : OAI22_X1 port map( A1 => n20448, A2 => n19716, B1 => n4819, B2 => 
                           n19727, ZN => n7758);
   U5400 : OAI22_X1 port map( A1 => n20451, A2 => n19716, B1 => n4818, B2 => 
                           n19726, ZN => n7759);
   U5401 : OAI22_X1 port map( A1 => n20454, A2 => n19716, B1 => n4817, B2 => 
                           n19726, ZN => n7760);
   U5402 : OAI22_X1 port map( A1 => n20457, A2 => n19716, B1 => n4816, B2 => 
                           n19726, ZN => n7761);
   U5403 : OAI22_X1 port map( A1 => n20460, A2 => n19716, B1 => n4815, B2 => 
                           n19726, ZN => n7762);
   U5404 : OAI22_X1 port map( A1 => n20463, A2 => n19716, B1 => n4814, B2 => 
                           n19725, ZN => n7763);
   U5405 : OAI22_X1 port map( A1 => n20466, A2 => n19716, B1 => n4813, B2 => 
                           n19725, ZN => n7764);
   U5406 : OAI22_X1 port map( A1 => n20469, A2 => n19716, B1 => n4812, B2 => 
                           n19725, ZN => n7765);
   U5407 : OAI22_X1 port map( A1 => n20472, A2 => n19716, B1 => n4811, B2 => 
                           n19725, ZN => n7766);
   U5408 : OAI22_X1 port map( A1 => n20475, A2 => n19718, B1 => n4810, B2 => 
                           n19724, ZN => n7767);
   U5409 : OAI22_X1 port map( A1 => n20478, A2 => n19717, B1 => n4809, B2 => 
                           n19724, ZN => n7768);
   U5410 : OAI22_X1 port map( A1 => n20481, A2 => n19716, B1 => n4808, B2 => 
                           n19724, ZN => n7769);
   U5411 : OAI22_X1 port map( A1 => n20484, A2 => n19718, B1 => n4807, B2 => 
                           n19724, ZN => n7770);
   U5412 : OAI22_X1 port map( A1 => n20487, A2 => n19717, B1 => n4806, B2 => 
                           n19723, ZN => n7771);
   U5413 : OAI22_X1 port map( A1 => n20490, A2 => n19716, B1 => n4805, B2 => 
                           n19723, ZN => n7772);
   U5414 : OAI22_X1 port map( A1 => n20493, A2 => n19718, B1 => n4804, B2 => 
                           n19723, ZN => n7773);
   U5415 : OAI22_X1 port map( A1 => n20496, A2 => n19717, B1 => n4803, B2 => 
                           n19723, ZN => n7774);
   U5416 : OAI22_X1 port map( A1 => n20499, A2 => n19716, B1 => n4802, B2 => 
                           n19722, ZN => n7775);
   U5417 : OAI22_X1 port map( A1 => n20502, A2 => n19718, B1 => n4801, B2 => 
                           n19722, ZN => n7776);
   U5418 : OAI22_X1 port map( A1 => n20505, A2 => n19717, B1 => n4800, B2 => 
                           n19722, ZN => n7777);
   U5419 : OAI22_X1 port map( A1 => n20508, A2 => n19717, B1 => n4799, B2 => 
                           n19722, ZN => n7778);
   U5420 : OAI22_X1 port map( A1 => n20511, A2 => n19718, B1 => n4798, B2 => 
                           n19721, ZN => n7779);
   U5421 : OAI22_X1 port map( A1 => n20514, A2 => n19717, B1 => n4797, B2 => 
                           n19721, ZN => n7780);
   U5422 : OAI22_X1 port map( A1 => n20517, A2 => n19716, B1 => n4796, B2 => 
                           n19721, ZN => n7781);
   U5423 : OAI22_X1 port map( A1 => n20520, A2 => n19716, B1 => n4795, B2 => 
                           n19721, ZN => n7782);
   U5424 : OAI22_X1 port map( A1 => n20523, A2 => n19718, B1 => n4794, B2 => 
                           n19720, ZN => n7783);
   U5425 : OAI22_X1 port map( A1 => n20526, A2 => n19717, B1 => n4793, B2 => 
                           n19720, ZN => n7784);
   U5426 : OAI22_X1 port map( A1 => n20529, A2 => n19716, B1 => n4792, B2 => 
                           n19720, ZN => n7785);
   U5427 : OAI22_X1 port map( A1 => n20532, A2 => n19718, B1 => n4791, B2 => 
                           n19720, ZN => n7786);
   U5428 : OAI22_X1 port map( A1 => n20535, A2 => n19718, B1 => n4790, B2 => 
                           n19719, ZN => n7787);
   U5429 : OAI22_X1 port map( A1 => n20538, A2 => n19717, B1 => n4789, B2 => 
                           n19719, ZN => n7788);
   U5430 : OAI22_X1 port map( A1 => n20541, A2 => n19716, B1 => n4788, B2 => 
                           n19719, ZN => n7789);
   U5431 : OAI22_X1 port map( A1 => n20572, A2 => n19717, B1 => n4787, B2 => 
                           n19719, ZN => n7790);
   U5432 : OAI22_X1 port map( A1 => n20355, A2 => n19717, B1 => n4850, B2 => 
                           n19734, ZN => n7727);
   U5433 : OAI22_X1 port map( A1 => n20358, A2 => n19716, B1 => n4849, B2 => 
                           n19734, ZN => n7728);
   U5434 : OAI22_X1 port map( A1 => n20361, A2 => n19716, B1 => n4848, B2 => 
                           n19734, ZN => n7729);
   U5435 : OAI22_X1 port map( A1 => n20364, A2 => n19718, B1 => n4847, B2 => 
                           n19734, ZN => n7730);
   U5436 : AOI22_X1 port map( A1 => n19231, A2 => registers_4_0_port, B1 => 
                           n19225, B2 => n11593, ZN => n11638);
   U5437 : AOI22_X1 port map( A1 => n19231, A2 => registers_4_1_port, B1 => 
                           n19225, B2 => n11501, ZN => n11525);
   U5438 : AOI22_X1 port map( A1 => n19231, A2 => registers_4_2_port, B1 => 
                           n19225, B2 => n11433, ZN => n11458);
   U5439 : AOI22_X1 port map( A1 => n19231, A2 => registers_4_3_port, B1 => 
                           n19225, B2 => n11366, ZN => n11391);
   U5440 : AOI22_X1 port map( A1 => n19231, A2 => registers_4_4_port, B1 => 
                           n19225, B2 => n17996, ZN => n11323);
   U5441 : AOI22_X1 port map( A1 => n19231, A2 => registers_4_5_port, B1 => 
                           n19225, B2 => n17997, ZN => n11256);
   U5442 : AOI22_X1 port map( A1 => n19231, A2 => registers_4_6_port, B1 => 
                           n19225, B2 => n17998, ZN => n11189);
   U5443 : AOI22_X1 port map( A1 => n19231, A2 => registers_4_7_port, B1 => 
                           n19225, B2 => n17999, ZN => n11122);
   U5444 : AOI22_X1 port map( A1 => n19231, A2 => registers_4_8_port, B1 => 
                           n19225, B2 => n18000, ZN => n11054);
   U5445 : AOI22_X1 port map( A1 => n19231, A2 => registers_4_9_port, B1 => 
                           n19225, B2 => n18001, ZN => n10987);
   U5446 : AOI22_X1 port map( A1 => n19231, A2 => registers_4_10_port, B1 => 
                           n19225, B2 => n18002, ZN => n10920);
   U5447 : AOI22_X1 port map( A1 => n19231, A2 => registers_4_11_port, B1 => 
                           n19225, B2 => n18003, ZN => n10852);
   U5448 : AOI22_X1 port map( A1 => n19232, A2 => registers_4_12_port, B1 => 
                           n19226, B2 => n18004, ZN => n10785);
   U5449 : AOI22_X1 port map( A1 => n19232, A2 => registers_4_13_port, B1 => 
                           n19226, B2 => n18005, ZN => n10718);
   U5450 : AOI22_X1 port map( A1 => n19232, A2 => registers_4_14_port, B1 => 
                           n19226, B2 => n18006, ZN => n10651);
   U5451 : AOI22_X1 port map( A1 => n19232, A2 => registers_4_15_port, B1 => 
                           n19226, B2 => n18007, ZN => n10583);
   U5452 : AOI22_X1 port map( A1 => n19232, A2 => registers_4_16_port, B1 => 
                           n19226, B2 => n18008, ZN => n10516);
   U5453 : AOI22_X1 port map( A1 => n19232, A2 => registers_4_17_port, B1 => 
                           n19226, B2 => n18009, ZN => n10449);
   U5454 : AOI22_X1 port map( A1 => n19232, A2 => registers_4_18_port, B1 => 
                           n19226, B2 => n18010, ZN => n10382);
   U5455 : AOI22_X1 port map( A1 => n19232, A2 => registers_4_19_port, B1 => 
                           n19226, B2 => n18011, ZN => n10314);
   U5456 : AOI22_X1 port map( A1 => n19232, A2 => registers_4_20_port, B1 => 
                           n19226, B2 => n18012, ZN => n10247);
   U5457 : AOI22_X1 port map( A1 => n19232, A2 => registers_4_21_port, B1 => 
                           n19226, B2 => n18013, ZN => n10180);
   U5458 : AOI22_X1 port map( A1 => n19232, A2 => registers_4_22_port, B1 => 
                           n19226, B2 => n18014, ZN => n10113);
   U5459 : AOI22_X1 port map( A1 => n19232, A2 => registers_4_23_port, B1 => 
                           n19226, B2 => n18015, ZN => n10045);
   U5460 : AOI22_X1 port map( A1 => n19233, A2 => registers_4_24_port, B1 => 
                           n19227, B2 => n18016, ZN => n9978);
   U5461 : AOI22_X1 port map( A1 => n19233, A2 => registers_4_25_port, B1 => 
                           n19227, B2 => n18017, ZN => n9911);
   U5462 : AOI22_X1 port map( A1 => n19233, A2 => registers_4_26_port, B1 => 
                           n19227, B2 => n18018, ZN => n9843);
   U5463 : AOI22_X1 port map( A1 => n19233, A2 => registers_4_27_port, B1 => 
                           n19227, B2 => n18019, ZN => n9776);
   U5464 : AOI22_X1 port map( A1 => n19233, A2 => registers_4_28_port, B1 => 
                           n19227, B2 => n18020, ZN => n9709);
   U5465 : AOI22_X1 port map( A1 => n19233, A2 => registers_4_29_port, B1 => 
                           n19227, B2 => n18021, ZN => n9642);
   U5466 : AOI22_X1 port map( A1 => n19233, A2 => registers_4_30_port, B1 => 
                           n19227, B2 => n18022, ZN => n9574);
   U5467 : AOI22_X1 port map( A1 => n19233, A2 => registers_4_31_port, B1 => 
                           n19227, B2 => n18023, ZN => n9507);
   U5468 : AOI22_X1 port map( A1 => n19233, A2 => registers_4_32_port, B1 => 
                           n19227, B2 => n18024, ZN => n9440);
   U5469 : AOI22_X1 port map( A1 => n19233, A2 => registers_4_33_port, B1 => 
                           n19227, B2 => n18025, ZN => n9373);
   U5470 : AOI22_X1 port map( A1 => n19233, A2 => registers_4_34_port, B1 => 
                           n19227, B2 => n18026, ZN => n9305);
   U5471 : AOI22_X1 port map( A1 => n19233, A2 => registers_4_35_port, B1 => 
                           n19227, B2 => n18027, ZN => n6998);
   U5472 : AOI22_X1 port map( A1 => n19234, A2 => registers_4_36_port, B1 => 
                           n19228, B2 => n18028, ZN => n6931);
   U5473 : AOI22_X1 port map( A1 => n19234, A2 => registers_4_37_port, B1 => 
                           n19228, B2 => n18029, ZN => n6864);
   U5474 : AOI22_X1 port map( A1 => n19234, A2 => registers_4_38_port, B1 => 
                           n19228, B2 => n18030, ZN => n6797);
   U5475 : AOI22_X1 port map( A1 => n19234, A2 => registers_4_39_port, B1 => 
                           n19228, B2 => n18031, ZN => n6730);
   U5476 : AOI22_X1 port map( A1 => n19234, A2 => registers_4_40_port, B1 => 
                           n19228, B2 => n18032, ZN => n6663);
   U5477 : AOI22_X1 port map( A1 => n19234, A2 => registers_4_41_port, B1 => 
                           n19228, B2 => n18033, ZN => n6596);
   U5478 : AOI22_X1 port map( A1 => n19234, A2 => registers_4_42_port, B1 => 
                           n19228, B2 => n18034, ZN => n6530);
   U5479 : AOI22_X1 port map( A1 => n19234, A2 => registers_4_43_port, B1 => 
                           n19228, B2 => n18035, ZN => n6464);
   U5480 : AOI22_X1 port map( A1 => n19234, A2 => registers_4_44_port, B1 => 
                           n19228, B2 => n18036, ZN => n6398);
   U5481 : AOI22_X1 port map( A1 => n19234, A2 => registers_4_45_port, B1 => 
                           n19228, B2 => n18037, ZN => n6332);
   U5482 : AOI22_X1 port map( A1 => n19234, A2 => registers_4_46_port, B1 => 
                           n19228, B2 => n18038, ZN => n6266);
   U5483 : AOI22_X1 port map( A1 => n19234, A2 => registers_4_47_port, B1 => 
                           n19228, B2 => n18039, ZN => n6200);
   U5484 : AOI22_X1 port map( A1 => n19235, A2 => registers_4_48_port, B1 => 
                           n19229, B2 => n18040, ZN => n6134);
   U5485 : AOI22_X1 port map( A1 => n19235, A2 => registers_4_49_port, B1 => 
                           n19229, B2 => n18041, ZN => n6068);
   U5486 : AOI22_X1 port map( A1 => n19235, A2 => registers_4_50_port, B1 => 
                           n19229, B2 => n18042, ZN => n6000);
   U5487 : AOI22_X1 port map( A1 => n19235, A2 => registers_4_51_port, B1 => 
                           n19229, B2 => n18043, ZN => n5932);
   U5488 : AOI22_X1 port map( A1 => n19235, A2 => registers_4_52_port, B1 => 
                           n19229, B2 => n18044, ZN => n5865);
   U5489 : AOI22_X1 port map( A1 => n19235, A2 => registers_4_53_port, B1 => 
                           n19229, B2 => n18045, ZN => n5798);
   U5490 : AOI22_X1 port map( A1 => n19235, A2 => registers_4_54_port, B1 => 
                           n19229, B2 => n18046, ZN => n5726);
   U5491 : AOI22_X1 port map( A1 => n19235, A2 => registers_4_55_port, B1 => 
                           n19229, B2 => n18047, ZN => n5656);
   U5492 : AOI22_X1 port map( A1 => n19235, A2 => registers_4_56_port, B1 => 
                           n19229, B2 => n18048, ZN => n5588);
   U5493 : AOI22_X1 port map( A1 => n19235, A2 => registers_4_57_port, B1 => 
                           n19229, B2 => n18049, ZN => n5519);
   U5494 : AOI22_X1 port map( A1 => n19235, A2 => registers_4_58_port, B1 => 
                           n19229, B2 => n18050, ZN => n5450);
   U5495 : AOI22_X1 port map( A1 => n19235, A2 => registers_4_59_port, B1 => 
                           n19229, B2 => n18051, ZN => n5382);
   U5496 : AOI22_X1 port map( A1 => n19236, A2 => registers_4_60_port, B1 => 
                           n19230, B2 => n18052, ZN => n5312);
   U5497 : AOI22_X1 port map( A1 => n19435, A2 => registers_4_60_port, B1 => 
                           n19429, B2 => n18052, ZN => n5188);
   U5498 : AOI22_X1 port map( A1 => n19236, A2 => registers_4_61_port, B1 => 
                           n19230, B2 => n18053, ZN => n4379);
   U5499 : AOI22_X1 port map( A1 => n19435, A2 => registers_4_61_port, B1 => 
                           n19429, B2 => n18053, ZN => n3906);
   U5500 : AOI22_X1 port map( A1 => n19236, A2 => registers_4_62_port, B1 => 
                           n19230, B2 => n18054, ZN => n3282);
   U5501 : AOI22_X1 port map( A1 => n19435, A2 => registers_4_62_port, B1 => 
                           n19429, B2 => n18054, ZN => n3232);
   U5502 : AOI22_X1 port map( A1 => n19236, A2 => registers_4_63_port, B1 => 
                           n19230, B2 => n18055, ZN => n3103);
   U5503 : AOI22_X1 port map( A1 => n19435, A2 => registers_4_63_port, B1 => 
                           n19429, B2 => n18055, ZN => n2981);
   U5504 : AOI22_X1 port map( A1 => n19017, A2 => registers_15_39_port, B1 => 
                           n19011, B2 => n6718, ZN => n6748);
   U5505 : AOI22_X1 port map( A1 => n19017, A2 => registers_15_40_port, B1 => 
                           n19011, B2 => n6651, ZN => n6681);
   U5506 : AOI22_X1 port map( A1 => n19017, A2 => registers_15_41_port, B1 => 
                           n19011, B2 => n6584, ZN => n6614);
   U5507 : AOI22_X1 port map( A1 => n19017, A2 => registers_15_42_port, B1 => 
                           n19011, B2 => n6518, ZN => n6548);
   U5508 : AOI22_X1 port map( A1 => n19017, A2 => registers_15_43_port, B1 => 
                           n19011, B2 => n6452, ZN => n6482);
   U5509 : AOI22_X1 port map( A1 => n19017, A2 => registers_15_44_port, B1 => 
                           n19011, B2 => n6386, ZN => n6416);
   U5510 : AOI22_X1 port map( A1 => n19017, A2 => registers_15_45_port, B1 => 
                           n19011, B2 => n6320, ZN => n6350);
   U5511 : AOI22_X1 port map( A1 => n19017, A2 => registers_15_46_port, B1 => 
                           n19011, B2 => n6254, ZN => n6284);
   U5512 : AOI22_X1 port map( A1 => n19017, A2 => registers_15_47_port, B1 => 
                           n19011, B2 => n6188, ZN => n6218);
   U5513 : AOI22_X1 port map( A1 => n19018, A2 => registers_15_48_port, B1 => 
                           n19012, B2 => n6122, ZN => n6152);
   U5514 : AOI22_X1 port map( A1 => n19018, A2 => registers_15_49_port, B1 => 
                           n19012, B2 => n6056, ZN => n6086);
   U5515 : AOI22_X1 port map( A1 => n19018, A2 => registers_15_50_port, B1 => 
                           n19012, B2 => n5988, ZN => n6018);
   U5516 : AOI22_X1 port map( A1 => n19018, A2 => registers_15_51_port, B1 => 
                           n19012, B2 => n5920, ZN => n5950);
   U5517 : AOI22_X1 port map( A1 => n19018, A2 => registers_15_52_port, B1 => 
                           n19012, B2 => n5853, ZN => n5883);
   U5518 : AOI22_X1 port map( A1 => n19018, A2 => registers_15_53_port, B1 => 
                           n19012, B2 => n5786, ZN => n5816);
   U5519 : AOI22_X1 port map( A1 => n19018, A2 => registers_15_54_port, B1 => 
                           n19012, B2 => n5714, ZN => n5744);
   U5520 : AOI22_X1 port map( A1 => n19018, A2 => registers_15_55_port, B1 => 
                           n19012, B2 => n5644, ZN => n5674);
   U5521 : AOI22_X1 port map( A1 => n19018, A2 => registers_15_56_port, B1 => 
                           n19012, B2 => n5576, ZN => n5606);
   U5522 : AOI22_X1 port map( A1 => n19018, A2 => registers_15_57_port, B1 => 
                           n19012, B2 => n5507, ZN => n5537);
   U5523 : AOI22_X1 port map( A1 => n19018, A2 => registers_15_58_port, B1 => 
                           n19012, B2 => n5438, ZN => n5468);
   U5524 : AOI22_X1 port map( A1 => n19018, A2 => registers_15_59_port, B1 => 
                           n19012, B2 => n5370, ZN => n5400);
   U5525 : AOI22_X1 port map( A1 => n19014, A2 => registers_15_0_port, B1 => 
                           n19008, B2 => n11618, ZN => n11685);
   U5526 : AOI22_X1 port map( A1 => n19014, A2 => registers_15_1_port, B1 => 
                           n19008, B2 => n11513, ZN => n11544);
   U5527 : AOI22_X1 port map( A1 => n19014, A2 => registers_15_2_port, B1 => 
                           n19008, B2 => n11446, ZN => n11476);
   U5528 : AOI22_X1 port map( A1 => n19014, A2 => registers_15_3_port, B1 => 
                           n19008, B2 => n11378, ZN => n11409);
   U5529 : AOI22_X1 port map( A1 => n19014, A2 => registers_15_4_port, B1 => 
                           n19008, B2 => n11311, ZN => n11342);
   U5530 : AOI22_X1 port map( A1 => n19014, A2 => registers_15_5_port, B1 => 
                           n19008, B2 => n11244, ZN => n11274);
   U5531 : AOI22_X1 port map( A1 => n19014, A2 => registers_15_6_port, B1 => 
                           n19008, B2 => n11177, ZN => n11207);
   U5532 : AOI22_X1 port map( A1 => n19014, A2 => registers_15_7_port, B1 => 
                           n19008, B2 => n11109, ZN => n11140);
   U5533 : AOI22_X1 port map( A1 => n19014, A2 => registers_15_8_port, B1 => 
                           n19008, B2 => n11042, ZN => n11073);
   U5534 : AOI22_X1 port map( A1 => n19014, A2 => registers_15_9_port, B1 => 
                           n19008, B2 => n10975, ZN => n11005);
   U5535 : AOI22_X1 port map( A1 => n19014, A2 => registers_15_10_port, B1 => 
                           n19008, B2 => n10908, ZN => n10938);
   U5536 : AOI22_X1 port map( A1 => n19014, A2 => registers_15_11_port, B1 => 
                           n19008, B2 => n10840, ZN => n10871);
   U5537 : AOI22_X1 port map( A1 => n19015, A2 => registers_15_12_port, B1 => 
                           n19009, B2 => n10773, ZN => n10804);
   U5538 : AOI22_X1 port map( A1 => n19015, A2 => registers_15_13_port, B1 => 
                           n19009, B2 => n10706, ZN => n10736);
   U5539 : AOI22_X1 port map( A1 => n19015, A2 => registers_15_14_port, B1 => 
                           n19009, B2 => n10638, ZN => n10669);
   U5540 : AOI22_X1 port map( A1 => n19015, A2 => registers_15_15_port, B1 => 
                           n19009, B2 => n10571, ZN => n10602);
   U5541 : AOI22_X1 port map( A1 => n19015, A2 => registers_15_16_port, B1 => 
                           n19009, B2 => n10504, ZN => n10534);
   U5542 : AOI22_X1 port map( A1 => n19015, A2 => registers_15_17_port, B1 => 
                           n19009, B2 => n10437, ZN => n10467);
   U5543 : AOI22_X1 port map( A1 => n19015, A2 => registers_15_18_port, B1 => 
                           n19009, B2 => n10369, ZN => n10400);
   U5544 : AOI22_X1 port map( A1 => n19015, A2 => registers_15_19_port, B1 => 
                           n19009, B2 => n10302, ZN => n10333);
   U5545 : AOI22_X1 port map( A1 => n19015, A2 => registers_15_20_port, B1 => 
                           n19009, B2 => n10235, ZN => n10265);
   U5546 : AOI22_X1 port map( A1 => n19015, A2 => registers_15_21_port, B1 => 
                           n19009, B2 => n10168, ZN => n10198);
   U5547 : AOI22_X1 port map( A1 => n19015, A2 => registers_15_22_port, B1 => 
                           n19009, B2 => n10100, ZN => n10131);
   U5548 : AOI22_X1 port map( A1 => n19015, A2 => registers_15_23_port, B1 => 
                           n19009, B2 => n10033, ZN => n10064);
   U5549 : AOI22_X1 port map( A1 => n19016, A2 => registers_15_24_port, B1 => 
                           n19010, B2 => n9966, ZN => n9996);
   U5550 : AOI22_X1 port map( A1 => n19016, A2 => registers_15_25_port, B1 => 
                           n19010, B2 => n9898, ZN => n9929);
   U5551 : AOI22_X1 port map( A1 => n19016, A2 => registers_15_26_port, B1 => 
                           n19010, B2 => n9831, ZN => n9862);
   U5552 : AOI22_X1 port map( A1 => n19016, A2 => registers_15_27_port, B1 => 
                           n19010, B2 => n9764, ZN => n9794);
   U5553 : AOI22_X1 port map( A1 => n19016, A2 => registers_15_28_port, B1 => 
                           n19010, B2 => n9697, ZN => n9727);
   U5554 : AOI22_X1 port map( A1 => n19016, A2 => registers_15_29_port, B1 => 
                           n19010, B2 => n9629, ZN => n9660);
   U5555 : AOI22_X1 port map( A1 => n19016, A2 => registers_15_30_port, B1 => 
                           n19010, B2 => n9562, ZN => n9593);
   U5556 : AOI22_X1 port map( A1 => n19016, A2 => registers_15_31_port, B1 => 
                           n19010, B2 => n9495, ZN => n9525);
   U5557 : AOI22_X1 port map( A1 => n19016, A2 => registers_15_32_port, B1 => 
                           n19010, B2 => n9428, ZN => n9458);
   U5558 : AOI22_X1 port map( A1 => n19016, A2 => registers_15_33_port, B1 => 
                           n19010, B2 => n9360, ZN => n9391);
   U5559 : AOI22_X1 port map( A1 => n19016, A2 => registers_15_34_port, B1 => 
                           n19010, B2 => n9293, ZN => n9324);
   U5560 : AOI22_X1 port map( A1 => n19016, A2 => registers_15_35_port, B1 => 
                           n19010, B2 => n6986, ZN => n7016);
   U5561 : AOI22_X1 port map( A1 => n19019, A2 => registers_15_60_port, B1 => 
                           n19013, B2 => n5300, ZN => n5330);
   U5562 : AOI22_X1 port map( A1 => n19019, A2 => registers_15_61_port, B1 => 
                           n19013, B2 => n4175, ZN => n4653);
   U5563 : AOI22_X1 port map( A1 => n19019, A2 => registers_15_62_port, B1 => 
                           n19013, B2 => n3258, ZN => n3435);
   U5564 : AOI22_X1 port map( A1 => n19019, A2 => registers_15_63_port, B1 => 
                           n19013, B2 => n3018, ZN => n3157);
   U5565 : AOI22_X1 port map( A1 => n19017, A2 => registers_15_36_port, B1 => 
                           n19011, B2 => n6919, ZN => n6950);
   U5566 : AOI22_X1 port map( A1 => n19017, A2 => registers_15_37_port, B1 => 
                           n19011, B2 => n6852, ZN => n6883);
   U5567 : OAI22_X1 port map( A1 => n20469, A2 => n19521, B1 => n5282, B2 => 
                           n19529, ZN => n7317);
   U5568 : OAI22_X1 port map( A1 => n20369, A2 => n20334, B1 => n3362, B2 => 
                           n20349, ZN => n9139);
   U5569 : OAI22_X1 port map( A1 => n20372, A2 => n20334, B1 => n3361, B2 => 
                           n20349, ZN => n9140);
   U5570 : OAI22_X1 port map( A1 => n20375, A2 => n20334, B1 => n3360, B2 => 
                           n20349, ZN => n9141);
   U5571 : OAI22_X1 port map( A1 => n20378, A2 => n20334, B1 => n3359, B2 => 
                           n20349, ZN => n9142);
   U5572 : OAI22_X1 port map( A1 => n20381, A2 => n20334, B1 => n3358, B2 => 
                           n20348, ZN => n9143);
   U5573 : OAI22_X1 port map( A1 => n20384, A2 => n20334, B1 => n3357, B2 => 
                           n20348, ZN => n9144);
   U5574 : OAI22_X1 port map( A1 => n20387, A2 => n20334, B1 => n3356, B2 => 
                           n20348, ZN => n9145);
   U5575 : OAI22_X1 port map( A1 => n20390, A2 => n20334, B1 => n3355, B2 => 
                           n20348, ZN => n9146);
   U5576 : OAI22_X1 port map( A1 => n20393, A2 => n20334, B1 => n3354, B2 => 
                           n20347, ZN => n9147);
   U5577 : OAI22_X1 port map( A1 => n20396, A2 => n20334, B1 => n3353, B2 => 
                           n20347, ZN => n9148);
   U5578 : OAI22_X1 port map( A1 => n20399, A2 => n20334, B1 => n3352, B2 => 
                           n20347, ZN => n9149);
   U5579 : OAI22_X1 port map( A1 => n20402, A2 => n20334, B1 => n3351, B2 => 
                           n20347, ZN => n9150);
   U5580 : OAI22_X1 port map( A1 => n20405, A2 => n20333, B1 => n3350, B2 => 
                           n20346, ZN => n9151);
   U5581 : OAI22_X1 port map( A1 => n20408, A2 => n20333, B1 => n3349, B2 => 
                           n20346, ZN => n9152);
   U5582 : OAI22_X1 port map( A1 => n20411, A2 => n20333, B1 => n3348, B2 => 
                           n20346, ZN => n9153);
   U5583 : OAI22_X1 port map( A1 => n20414, A2 => n20333, B1 => n3347, B2 => 
                           n20346, ZN => n9154);
   U5584 : OAI22_X1 port map( A1 => n20417, A2 => n20333, B1 => n3346, B2 => 
                           n20345, ZN => n9155);
   U5585 : OAI22_X1 port map( A1 => n20420, A2 => n20333, B1 => n3345, B2 => 
                           n20345, ZN => n9156);
   U5586 : OAI22_X1 port map( A1 => n20423, A2 => n20333, B1 => n3344, B2 => 
                           n20345, ZN => n9157);
   U5587 : OAI22_X1 port map( A1 => n20426, A2 => n20333, B1 => n3343, B2 => 
                           n20345, ZN => n9158);
   U5588 : OAI22_X1 port map( A1 => n20429, A2 => n20333, B1 => n3342, B2 => 
                           n20344, ZN => n9159);
   U5589 : OAI22_X1 port map( A1 => n20432, A2 => n20333, B1 => n3341, B2 => 
                           n20344, ZN => n9160);
   U5590 : OAI22_X1 port map( A1 => n20435, A2 => n20333, B1 => n3340, B2 => 
                           n20344, ZN => n9161);
   U5591 : OAI22_X1 port map( A1 => n20438, A2 => n20333, B1 => n3339, B2 => 
                           n20344, ZN => n9162);
   U5592 : OAI22_X1 port map( A1 => n20441, A2 => n20332, B1 => n3338, B2 => 
                           n20343, ZN => n9163);
   U5593 : OAI22_X1 port map( A1 => n20444, A2 => n20332, B1 => n3337, B2 => 
                           n20343, ZN => n9164);
   U5594 : OAI22_X1 port map( A1 => n20447, A2 => n20332, B1 => n3336, B2 => 
                           n20343, ZN => n9165);
   U5595 : OAI22_X1 port map( A1 => n20450, A2 => n20332, B1 => n3335, B2 => 
                           n20343, ZN => n9166);
   U5596 : OAI22_X1 port map( A1 => n20453, A2 => n20332, B1 => n3334, B2 => 
                           n20342, ZN => n9167);
   U5597 : OAI22_X1 port map( A1 => n20456, A2 => n20332, B1 => n3333, B2 => 
                           n20342, ZN => n9168);
   U5598 : OAI22_X1 port map( A1 => n20459, A2 => n20332, B1 => n3332, B2 => 
                           n20342, ZN => n9169);
   U5599 : OAI22_X1 port map( A1 => n20462, A2 => n20332, B1 => n3331, B2 => 
                           n20342, ZN => n9170);
   U5600 : OAI22_X1 port map( A1 => n20465, A2 => n20332, B1 => n3330, B2 => 
                           n20341, ZN => n9171);
   U5601 : OAI22_X1 port map( A1 => n20468, A2 => n20332, B1 => n3329, B2 => 
                           n20341, ZN => n9172);
   U5602 : OAI22_X1 port map( A1 => n20471, A2 => n20332, B1 => n3328, B2 => 
                           n20341, ZN => n9173);
   U5603 : OAI22_X1 port map( A1 => n20474, A2 => n20332, B1 => n3327, B2 => 
                           n20341, ZN => n9174);
   U5604 : OAI22_X1 port map( A1 => n20477, A2 => n20334, B1 => n3326, B2 => 
                           n20340, ZN => n9175);
   U5605 : OAI22_X1 port map( A1 => n20480, A2 => n20333, B1 => n3325, B2 => 
                           n20340, ZN => n9176);
   U5606 : OAI22_X1 port map( A1 => n20483, A2 => n20332, B1 => n3324, B2 => 
                           n20340, ZN => n9177);
   U5607 : OAI22_X1 port map( A1 => n20486, A2 => n20332, B1 => n3323, B2 => 
                           n20340, ZN => n9178);
   U5608 : OAI22_X1 port map( A1 => n20489, A2 => n20334, B1 => n3322, B2 => 
                           n20339, ZN => n9179);
   U5609 : OAI22_X1 port map( A1 => n20492, A2 => n20333, B1 => n3321, B2 => 
                           n20339, ZN => n9180);
   U5610 : OAI22_X1 port map( A1 => n20495, A2 => n20332, B1 => n3320, B2 => 
                           n20339, ZN => n9181);
   U5611 : OAI22_X1 port map( A1 => n20498, A2 => n20334, B1 => n3319, B2 => 
                           n20339, ZN => n9182);
   U5612 : OAI22_X1 port map( A1 => n20501, A2 => n20334, B1 => n3318, B2 => 
                           n20338, ZN => n9183);
   U5613 : OAI22_X1 port map( A1 => n20504, A2 => n20333, B1 => n3317, B2 => 
                           n20338, ZN => n9184);
   U5614 : OAI22_X1 port map( A1 => n20507, A2 => n20332, B1 => n3316, B2 => 
                           n20338, ZN => n9185);
   U5615 : OAI22_X1 port map( A1 => n20510, A2 => n20333, B1 => n3315, B2 => 
                           n20338, ZN => n9186);
   U5616 : OAI22_X1 port map( A1 => n20513, A2 => n20334, B1 => n3314, B2 => 
                           n20337, ZN => n9187);
   U5617 : OAI22_X1 port map( A1 => n20516, A2 => n20333, B1 => n3313, B2 => 
                           n20337, ZN => n9188);
   U5618 : OAI22_X1 port map( A1 => n20519, A2 => n20332, B1 => n3312, B2 => 
                           n20337, ZN => n9189);
   U5619 : OAI22_X1 port map( A1 => n20522, A2 => n20334, B1 => n3311, B2 => 
                           n20337, ZN => n9190);
   U5620 : OAI22_X1 port map( A1 => n20525, A2 => n20333, B1 => n3310, B2 => 
                           n20336, ZN => n9191);
   U5621 : OAI22_X1 port map( A1 => n20528, A2 => n20332, B1 => n3309, B2 => 
                           n20336, ZN => n9192);
   U5622 : OAI22_X1 port map( A1 => n20531, A2 => n20334, B1 => n3308, B2 => 
                           n20336, ZN => n9193);
   U5623 : OAI22_X1 port map( A1 => n20534, A2 => n20333, B1 => n3307, B2 => 
                           n20336, ZN => n9194);
   U5624 : OAI22_X1 port map( A1 => n20537, A2 => n20332, B1 => n3306, B2 => 
                           n20335, ZN => n9195);
   U5625 : OAI22_X1 port map( A1 => n20540, A2 => n20334, B1 => n3305, B2 => 
                           n20335, ZN => n9196);
   U5626 : OAI22_X1 port map( A1 => n20543, A2 => n20333, B1 => n3304, B2 => 
                           n20335, ZN => n9197);
   U5627 : OAI22_X1 port map( A1 => n20574, A2 => n20333, B1 => n3303, B2 => 
                           n20335, ZN => n9198);
   U5628 : OAI22_X1 port map( A1 => n20357, A2 => n20333, B1 => n3366, B2 => 
                           n20350, ZN => n9135);
   U5629 : OAI22_X1 port map( A1 => n20360, A2 => n20332, B1 => n3365, B2 => 
                           n20350, ZN => n9136);
   U5630 : OAI22_X1 port map( A1 => n20363, A2 => n20332, B1 => n3364, B2 => 
                           n20350, ZN => n9137);
   U5631 : OAI22_X1 port map( A1 => n20366, A2 => n20334, B1 => n3363, B2 => 
                           n20350, ZN => n9138);
   U5632 : OAI22_X1 port map( A1 => n20369, A2 => n20306, B1 => n3430, B2 => 
                           n20321, ZN => n9075);
   U5633 : OAI22_X1 port map( A1 => n20372, A2 => n20306, B1 => n3429, B2 => 
                           n20321, ZN => n9076);
   U5634 : OAI22_X1 port map( A1 => n20375, A2 => n20306, B1 => n3428, B2 => 
                           n20321, ZN => n9077);
   U5635 : OAI22_X1 port map( A1 => n20378, A2 => n20306, B1 => n3427, B2 => 
                           n20321, ZN => n9078);
   U5636 : OAI22_X1 port map( A1 => n20381, A2 => n20306, B1 => n3426, B2 => 
                           n20320, ZN => n9079);
   U5637 : OAI22_X1 port map( A1 => n20384, A2 => n20306, B1 => n3425, B2 => 
                           n20320, ZN => n9080);
   U5638 : OAI22_X1 port map( A1 => n20387, A2 => n20306, B1 => n3424, B2 => 
                           n20320, ZN => n9081);
   U5639 : OAI22_X1 port map( A1 => n20390, A2 => n20306, B1 => n3423, B2 => 
                           n20320, ZN => n9082);
   U5640 : OAI22_X1 port map( A1 => n20393, A2 => n20306, B1 => n3422, B2 => 
                           n20319, ZN => n9083);
   U5641 : OAI22_X1 port map( A1 => n20396, A2 => n20306, B1 => n3421, B2 => 
                           n20319, ZN => n9084);
   U5642 : OAI22_X1 port map( A1 => n20399, A2 => n20306, B1 => n3420, B2 => 
                           n20319, ZN => n9085);
   U5643 : OAI22_X1 port map( A1 => n20402, A2 => n20306, B1 => n3419, B2 => 
                           n20319, ZN => n9086);
   U5644 : OAI22_X1 port map( A1 => n20405, A2 => n20305, B1 => n3418, B2 => 
                           n20318, ZN => n9087);
   U5645 : OAI22_X1 port map( A1 => n20408, A2 => n20305, B1 => n3417, B2 => 
                           n20318, ZN => n9088);
   U5646 : OAI22_X1 port map( A1 => n20411, A2 => n20305, B1 => n3416, B2 => 
                           n20318, ZN => n9089);
   U5647 : OAI22_X1 port map( A1 => n20414, A2 => n20305, B1 => n3415, B2 => 
                           n20318, ZN => n9090);
   U5648 : OAI22_X1 port map( A1 => n20417, A2 => n20305, B1 => n3414, B2 => 
                           n20317, ZN => n9091);
   U5649 : OAI22_X1 port map( A1 => n20420, A2 => n20305, B1 => n3413, B2 => 
                           n20317, ZN => n9092);
   U5650 : OAI22_X1 port map( A1 => n20423, A2 => n20305, B1 => n3412, B2 => 
                           n20317, ZN => n9093);
   U5651 : OAI22_X1 port map( A1 => n20426, A2 => n20305, B1 => n3411, B2 => 
                           n20317, ZN => n9094);
   U5652 : OAI22_X1 port map( A1 => n20429, A2 => n20305, B1 => n3410, B2 => 
                           n20316, ZN => n9095);
   U5653 : OAI22_X1 port map( A1 => n20432, A2 => n20305, B1 => n3409, B2 => 
                           n20316, ZN => n9096);
   U5654 : OAI22_X1 port map( A1 => n20435, A2 => n20305, B1 => n3408, B2 => 
                           n20316, ZN => n9097);
   U5655 : OAI22_X1 port map( A1 => n20438, A2 => n20305, B1 => n3407, B2 => 
                           n20316, ZN => n9098);
   U5656 : OAI22_X1 port map( A1 => n20441, A2 => n20304, B1 => n3406, B2 => 
                           n20315, ZN => n9099);
   U5657 : OAI22_X1 port map( A1 => n20444, A2 => n20304, B1 => n3405, B2 => 
                           n20315, ZN => n9100);
   U5658 : OAI22_X1 port map( A1 => n20447, A2 => n20304, B1 => n3404, B2 => 
                           n20315, ZN => n9101);
   U5659 : OAI22_X1 port map( A1 => n20450, A2 => n20304, B1 => n3403, B2 => 
                           n20315, ZN => n9102);
   U5660 : OAI22_X1 port map( A1 => n20453, A2 => n20304, B1 => n3402, B2 => 
                           n20314, ZN => n9103);
   U5661 : OAI22_X1 port map( A1 => n20456, A2 => n20304, B1 => n3401, B2 => 
                           n20314, ZN => n9104);
   U5662 : OAI22_X1 port map( A1 => n20459, A2 => n20304, B1 => n3400, B2 => 
                           n20314, ZN => n9105);
   U5663 : OAI22_X1 port map( A1 => n20462, A2 => n20304, B1 => n3399, B2 => 
                           n20314, ZN => n9106);
   U5664 : OAI22_X1 port map( A1 => n20465, A2 => n20304, B1 => n3398, B2 => 
                           n20313, ZN => n9107);
   U5665 : OAI22_X1 port map( A1 => n20468, A2 => n20304, B1 => n3397, B2 => 
                           n20313, ZN => n9108);
   U5666 : OAI22_X1 port map( A1 => n20471, A2 => n20304, B1 => n3396, B2 => 
                           n20313, ZN => n9109);
   U5667 : OAI22_X1 port map( A1 => n20474, A2 => n20304, B1 => n3395, B2 => 
                           n20313, ZN => n9110);
   U5668 : OAI22_X1 port map( A1 => n20477, A2 => n20306, B1 => n3394, B2 => 
                           n20312, ZN => n9111);
   U5669 : OAI22_X1 port map( A1 => n20480, A2 => n20305, B1 => n3393, B2 => 
                           n20312, ZN => n9112);
   U5670 : OAI22_X1 port map( A1 => n20483, A2 => n20304, B1 => n3392, B2 => 
                           n20312, ZN => n9113);
   U5671 : OAI22_X1 port map( A1 => n20486, A2 => n20306, B1 => n3391, B2 => 
                           n20312, ZN => n9114);
   U5672 : OAI22_X1 port map( A1 => n20489, A2 => n20305, B1 => n3390, B2 => 
                           n20311, ZN => n9115);
   U5673 : OAI22_X1 port map( A1 => n20492, A2 => n20304, B1 => n3389, B2 => 
                           n20311, ZN => n9116);
   U5674 : OAI22_X1 port map( A1 => n20495, A2 => n20306, B1 => n3388, B2 => 
                           n20311, ZN => n9117);
   U5675 : OAI22_X1 port map( A1 => n20498, A2 => n20305, B1 => n3387, B2 => 
                           n20311, ZN => n9118);
   U5676 : OAI22_X1 port map( A1 => n20501, A2 => n20304, B1 => n3386, B2 => 
                           n20310, ZN => n9119);
   U5677 : OAI22_X1 port map( A1 => n20504, A2 => n20306, B1 => n3385, B2 => 
                           n20310, ZN => n9120);
   U5678 : OAI22_X1 port map( A1 => n20507, A2 => n20305, B1 => n3384, B2 => 
                           n20310, ZN => n9121);
   U5679 : OAI22_X1 port map( A1 => n20510, A2 => n20305, B1 => n3383, B2 => 
                           n20310, ZN => n9122);
   U5680 : OAI22_X1 port map( A1 => n20513, A2 => n20306, B1 => n3382, B2 => 
                           n20309, ZN => n9123);
   U5681 : OAI22_X1 port map( A1 => n20516, A2 => n20305, B1 => n3381, B2 => 
                           n20309, ZN => n9124);
   U5682 : OAI22_X1 port map( A1 => n20519, A2 => n20304, B1 => n3380, B2 => 
                           n20309, ZN => n9125);
   U5683 : OAI22_X1 port map( A1 => n20522, A2 => n20304, B1 => n3379, B2 => 
                           n20309, ZN => n9126);
   U5684 : OAI22_X1 port map( A1 => n20525, A2 => n20306, B1 => n3378, B2 => 
                           n20308, ZN => n9127);
   U5685 : OAI22_X1 port map( A1 => n20528, A2 => n20305, B1 => n3377, B2 => 
                           n20308, ZN => n9128);
   U5686 : OAI22_X1 port map( A1 => n20531, A2 => n20304, B1 => n3376, B2 => 
                           n20308, ZN => n9129);
   U5687 : OAI22_X1 port map( A1 => n20534, A2 => n20306, B1 => n3375, B2 => 
                           n20308, ZN => n9130);
   U5688 : OAI22_X1 port map( A1 => n20537, A2 => n20306, B1 => n3374, B2 => 
                           n20307, ZN => n9131);
   U5689 : OAI22_X1 port map( A1 => n20540, A2 => n20305, B1 => n3373, B2 => 
                           n20307, ZN => n9132);
   U5690 : OAI22_X1 port map( A1 => n20543, A2 => n20304, B1 => n3372, B2 => 
                           n20307, ZN => n9133);
   U5691 : OAI22_X1 port map( A1 => n20574, A2 => n20305, B1 => n3371, B2 => 
                           n20307, ZN => n9134);
   U5692 : OAI22_X1 port map( A1 => n20357, A2 => n20305, B1 => n3434, B2 => 
                           n20322, ZN => n9071);
   U5693 : OAI22_X1 port map( A1 => n20360, A2 => n20304, B1 => n3433, B2 => 
                           n20322, ZN => n9072);
   U5694 : OAI22_X1 port map( A1 => n20363, A2 => n20304, B1 => n3432, B2 => 
                           n20322, ZN => n9073);
   U5695 : OAI22_X1 port map( A1 => n20366, A2 => n20306, B1 => n3431, B2 => 
                           n20322, ZN => n9074);
   U5696 : OAI22_X1 port map( A1 => n20369, A2 => n20166, B1 => n3766, B2 => 
                           n20181, ZN => n8755);
   U5697 : OAI22_X1 port map( A1 => n20372, A2 => n20166, B1 => n3765, B2 => 
                           n20181, ZN => n8756);
   U5698 : OAI22_X1 port map( A1 => n20375, A2 => n20166, B1 => n3764, B2 => 
                           n20181, ZN => n8757);
   U5699 : OAI22_X1 port map( A1 => n20378, A2 => n20166, B1 => n3763, B2 => 
                           n20181, ZN => n8758);
   U5700 : OAI22_X1 port map( A1 => n20381, A2 => n20166, B1 => n3762, B2 => 
                           n20180, ZN => n8759);
   U5701 : OAI22_X1 port map( A1 => n20384, A2 => n20166, B1 => n3761, B2 => 
                           n20180, ZN => n8760);
   U5702 : OAI22_X1 port map( A1 => n20387, A2 => n20166, B1 => n3760, B2 => 
                           n20180, ZN => n8761);
   U5703 : OAI22_X1 port map( A1 => n20390, A2 => n20166, B1 => n3759, B2 => 
                           n20180, ZN => n8762);
   U5704 : OAI22_X1 port map( A1 => n20393, A2 => n20166, B1 => n3758, B2 => 
                           n20179, ZN => n8763);
   U5705 : OAI22_X1 port map( A1 => n20396, A2 => n20166, B1 => n3757, B2 => 
                           n20179, ZN => n8764);
   U5706 : OAI22_X1 port map( A1 => n20399, A2 => n20166, B1 => n3756, B2 => 
                           n20179, ZN => n8765);
   U5707 : OAI22_X1 port map( A1 => n20402, A2 => n20166, B1 => n3755, B2 => 
                           n20179, ZN => n8766);
   U5708 : OAI22_X1 port map( A1 => n20405, A2 => n20165, B1 => n3754, B2 => 
                           n20178, ZN => n8767);
   U5709 : OAI22_X1 port map( A1 => n20408, A2 => n20165, B1 => n3753, B2 => 
                           n20178, ZN => n8768);
   U5710 : OAI22_X1 port map( A1 => n20411, A2 => n20165, B1 => n3752, B2 => 
                           n20178, ZN => n8769);
   U5711 : OAI22_X1 port map( A1 => n20414, A2 => n20165, B1 => n3751, B2 => 
                           n20178, ZN => n8770);
   U5712 : OAI22_X1 port map( A1 => n20417, A2 => n20165, B1 => n3750, B2 => 
                           n20177, ZN => n8771);
   U5713 : OAI22_X1 port map( A1 => n20420, A2 => n20165, B1 => n3749, B2 => 
                           n20177, ZN => n8772);
   U5714 : OAI22_X1 port map( A1 => n20423, A2 => n20165, B1 => n3748, B2 => 
                           n20177, ZN => n8773);
   U5715 : OAI22_X1 port map( A1 => n20426, A2 => n20165, B1 => n3747, B2 => 
                           n20177, ZN => n8774);
   U5716 : OAI22_X1 port map( A1 => n20429, A2 => n20165, B1 => n3746, B2 => 
                           n20176, ZN => n8775);
   U5717 : OAI22_X1 port map( A1 => n20432, A2 => n20165, B1 => n3745, B2 => 
                           n20176, ZN => n8776);
   U5718 : OAI22_X1 port map( A1 => n20435, A2 => n20165, B1 => n3744, B2 => 
                           n20176, ZN => n8777);
   U5719 : OAI22_X1 port map( A1 => n20438, A2 => n20165, B1 => n3743, B2 => 
                           n20176, ZN => n8778);
   U5720 : OAI22_X1 port map( A1 => n20441, A2 => n20164, B1 => n3742, B2 => 
                           n20175, ZN => n8779);
   U5721 : OAI22_X1 port map( A1 => n20444, A2 => n20164, B1 => n3741, B2 => 
                           n20175, ZN => n8780);
   U5722 : OAI22_X1 port map( A1 => n20447, A2 => n20164, B1 => n3740, B2 => 
                           n20175, ZN => n8781);
   U5723 : OAI22_X1 port map( A1 => n20450, A2 => n20164, B1 => n3739, B2 => 
                           n20175, ZN => n8782);
   U5724 : OAI22_X1 port map( A1 => n20453, A2 => n20164, B1 => n3738, B2 => 
                           n20174, ZN => n8783);
   U5725 : OAI22_X1 port map( A1 => n20456, A2 => n20164, B1 => n3737, B2 => 
                           n20174, ZN => n8784);
   U5726 : OAI22_X1 port map( A1 => n20459, A2 => n20164, B1 => n3736, B2 => 
                           n20174, ZN => n8785);
   U5727 : OAI22_X1 port map( A1 => n20462, A2 => n20164, B1 => n3735, B2 => 
                           n20174, ZN => n8786);
   U5728 : OAI22_X1 port map( A1 => n20465, A2 => n20164, B1 => n3734, B2 => 
                           n20173, ZN => n8787);
   U5729 : OAI22_X1 port map( A1 => n20468, A2 => n20164, B1 => n3733, B2 => 
                           n20173, ZN => n8788);
   U5730 : OAI22_X1 port map( A1 => n20471, A2 => n20164, B1 => n3732, B2 => 
                           n20173, ZN => n8789);
   U5731 : OAI22_X1 port map( A1 => n20474, A2 => n20164, B1 => n3731, B2 => 
                           n20173, ZN => n8790);
   U5732 : OAI22_X1 port map( A1 => n20477, A2 => n20166, B1 => n3730, B2 => 
                           n20172, ZN => n8791);
   U5733 : OAI22_X1 port map( A1 => n20480, A2 => n20165, B1 => n3729, B2 => 
                           n20172, ZN => n8792);
   U5734 : OAI22_X1 port map( A1 => n20483, A2 => n20164, B1 => n3728, B2 => 
                           n20172, ZN => n8793);
   U5735 : OAI22_X1 port map( A1 => n20486, A2 => n20166, B1 => n3727, B2 => 
                           n20172, ZN => n8794);
   U5736 : OAI22_X1 port map( A1 => n20489, A2 => n20165, B1 => n3726, B2 => 
                           n20171, ZN => n8795);
   U5737 : OAI22_X1 port map( A1 => n20492, A2 => n20164, B1 => n3725, B2 => 
                           n20171, ZN => n8796);
   U5738 : OAI22_X1 port map( A1 => n20495, A2 => n20166, B1 => n3724, B2 => 
                           n20171, ZN => n8797);
   U5739 : OAI22_X1 port map( A1 => n20498, A2 => n20165, B1 => n3723, B2 => 
                           n20171, ZN => n8798);
   U5740 : OAI22_X1 port map( A1 => n20501, A2 => n20164, B1 => n3722, B2 => 
                           n20170, ZN => n8799);
   U5741 : OAI22_X1 port map( A1 => n20504, A2 => n20166, B1 => n3721, B2 => 
                           n20170, ZN => n8800);
   U5742 : OAI22_X1 port map( A1 => n20507, A2 => n20165, B1 => n3720, B2 => 
                           n20170, ZN => n8801);
   U5743 : OAI22_X1 port map( A1 => n20510, A2 => n20165, B1 => n3719, B2 => 
                           n20170, ZN => n8802);
   U5744 : OAI22_X1 port map( A1 => n20513, A2 => n20166, B1 => n3718, B2 => 
                           n20169, ZN => n8803);
   U5745 : OAI22_X1 port map( A1 => n20516, A2 => n20165, B1 => n3717, B2 => 
                           n20169, ZN => n8804);
   U5746 : OAI22_X1 port map( A1 => n20519, A2 => n20164, B1 => n3716, B2 => 
                           n20169, ZN => n8805);
   U5747 : OAI22_X1 port map( A1 => n20522, A2 => n20164, B1 => n3715, B2 => 
                           n20169, ZN => n8806);
   U5748 : OAI22_X1 port map( A1 => n20525, A2 => n20166, B1 => n3714, B2 => 
                           n20168, ZN => n8807);
   U5749 : OAI22_X1 port map( A1 => n20528, A2 => n20165, B1 => n3713, B2 => 
                           n20168, ZN => n8808);
   U5750 : OAI22_X1 port map( A1 => n20531, A2 => n20164, B1 => n3712, B2 => 
                           n20168, ZN => n8809);
   U5751 : OAI22_X1 port map( A1 => n20534, A2 => n20166, B1 => n3711, B2 => 
                           n20168, ZN => n8810);
   U5752 : OAI22_X1 port map( A1 => n20537, A2 => n20166, B1 => n3710, B2 => 
                           n20167, ZN => n8811);
   U5753 : OAI22_X1 port map( A1 => n20540, A2 => n20165, B1 => n3709, B2 => 
                           n20167, ZN => n8812);
   U5754 : OAI22_X1 port map( A1 => n20543, A2 => n20164, B1 => n3708, B2 => 
                           n20167, ZN => n8813);
   U5755 : OAI22_X1 port map( A1 => n20574, A2 => n20165, B1 => n3707, B2 => 
                           n20167, ZN => n8814);
   U5756 : OAI22_X1 port map( A1 => n20357, A2 => n20165, B1 => n3770, B2 => 
                           n20182, ZN => n8751);
   U5757 : OAI22_X1 port map( A1 => n20360, A2 => n20164, B1 => n3769, B2 => 
                           n20182, ZN => n8752);
   U5758 : OAI22_X1 port map( A1 => n20363, A2 => n20164, B1 => n3768, B2 => 
                           n20182, ZN => n8753);
   U5759 : OAI22_X1 port map( A1 => n20366, A2 => n20166, B1 => n3767, B2 => 
                           n20182, ZN => n8754);
   U5760 : OAI22_X1 port map( A1 => n20369, A2 => n20278, B1 => n3498, B2 => 
                           n20293, ZN => n9011);
   U5761 : OAI22_X1 port map( A1 => n20372, A2 => n20278, B1 => n3497, B2 => 
                           n20293, ZN => n9012);
   U5762 : OAI22_X1 port map( A1 => n20375, A2 => n20278, B1 => n3496, B2 => 
                           n20293, ZN => n9013);
   U5763 : OAI22_X1 port map( A1 => n20378, A2 => n20278, B1 => n3495, B2 => 
                           n20293, ZN => n9014);
   U5764 : OAI22_X1 port map( A1 => n20381, A2 => n20278, B1 => n3494, B2 => 
                           n20292, ZN => n9015);
   U5765 : OAI22_X1 port map( A1 => n20384, A2 => n20278, B1 => n3493, B2 => 
                           n20292, ZN => n9016);
   U5766 : OAI22_X1 port map( A1 => n20387, A2 => n20278, B1 => n3492, B2 => 
                           n20292, ZN => n9017);
   U5767 : OAI22_X1 port map( A1 => n20390, A2 => n20278, B1 => n3491, B2 => 
                           n20292, ZN => n9018);
   U5768 : OAI22_X1 port map( A1 => n20393, A2 => n20278, B1 => n3490, B2 => 
                           n20291, ZN => n9019);
   U5769 : OAI22_X1 port map( A1 => n20396, A2 => n20278, B1 => n3489, B2 => 
                           n20291, ZN => n9020);
   U5770 : OAI22_X1 port map( A1 => n20399, A2 => n20278, B1 => n3488, B2 => 
                           n20291, ZN => n9021);
   U5771 : OAI22_X1 port map( A1 => n20402, A2 => n20278, B1 => n3487, B2 => 
                           n20291, ZN => n9022);
   U5772 : OAI22_X1 port map( A1 => n20405, A2 => n20277, B1 => n3486, B2 => 
                           n20290, ZN => n9023);
   U5773 : OAI22_X1 port map( A1 => n20408, A2 => n20277, B1 => n3485, B2 => 
                           n20290, ZN => n9024);
   U5774 : OAI22_X1 port map( A1 => n20411, A2 => n20277, B1 => n3484, B2 => 
                           n20290, ZN => n9025);
   U5775 : OAI22_X1 port map( A1 => n20414, A2 => n20277, B1 => n3483, B2 => 
                           n20290, ZN => n9026);
   U5776 : OAI22_X1 port map( A1 => n20417, A2 => n20277, B1 => n3482, B2 => 
                           n20289, ZN => n9027);
   U5777 : OAI22_X1 port map( A1 => n20420, A2 => n20277, B1 => n3481, B2 => 
                           n20289, ZN => n9028);
   U5778 : OAI22_X1 port map( A1 => n20423, A2 => n20277, B1 => n3480, B2 => 
                           n20289, ZN => n9029);
   U5779 : OAI22_X1 port map( A1 => n20426, A2 => n20277, B1 => n3479, B2 => 
                           n20289, ZN => n9030);
   U5780 : OAI22_X1 port map( A1 => n20429, A2 => n20277, B1 => n3478, B2 => 
                           n20288, ZN => n9031);
   U5781 : OAI22_X1 port map( A1 => n20432, A2 => n20277, B1 => n3477, B2 => 
                           n20288, ZN => n9032);
   U5782 : OAI22_X1 port map( A1 => n20435, A2 => n20277, B1 => n3476, B2 => 
                           n20288, ZN => n9033);
   U5783 : OAI22_X1 port map( A1 => n20438, A2 => n20277, B1 => n3475, B2 => 
                           n20288, ZN => n9034);
   U5784 : OAI22_X1 port map( A1 => n20441, A2 => n20276, B1 => n3474, B2 => 
                           n20287, ZN => n9035);
   U5785 : OAI22_X1 port map( A1 => n20444, A2 => n20276, B1 => n3473, B2 => 
                           n20287, ZN => n9036);
   U5786 : OAI22_X1 port map( A1 => n20447, A2 => n20276, B1 => n3472, B2 => 
                           n20287, ZN => n9037);
   U5787 : OAI22_X1 port map( A1 => n20450, A2 => n20276, B1 => n3471, B2 => 
                           n20287, ZN => n9038);
   U5788 : OAI22_X1 port map( A1 => n20453, A2 => n20276, B1 => n3470, B2 => 
                           n20286, ZN => n9039);
   U5789 : OAI22_X1 port map( A1 => n20456, A2 => n20276, B1 => n3469, B2 => 
                           n20286, ZN => n9040);
   U5790 : OAI22_X1 port map( A1 => n20459, A2 => n20276, B1 => n3468, B2 => 
                           n20286, ZN => n9041);
   U5791 : OAI22_X1 port map( A1 => n20462, A2 => n20276, B1 => n3467, B2 => 
                           n20286, ZN => n9042);
   U5792 : OAI22_X1 port map( A1 => n20465, A2 => n20276, B1 => n3466, B2 => 
                           n20285, ZN => n9043);
   U5793 : OAI22_X1 port map( A1 => n20468, A2 => n20276, B1 => n3465, B2 => 
                           n20285, ZN => n9044);
   U5794 : OAI22_X1 port map( A1 => n20471, A2 => n20276, B1 => n3464, B2 => 
                           n20285, ZN => n9045);
   U5795 : OAI22_X1 port map( A1 => n20474, A2 => n20276, B1 => n3463, B2 => 
                           n20285, ZN => n9046);
   U5796 : OAI22_X1 port map( A1 => n20477, A2 => n20278, B1 => n3462, B2 => 
                           n20284, ZN => n9047);
   U5797 : OAI22_X1 port map( A1 => n20480, A2 => n20277, B1 => n3461, B2 => 
                           n20284, ZN => n9048);
   U5798 : OAI22_X1 port map( A1 => n20483, A2 => n20276, B1 => n3460, B2 => 
                           n20284, ZN => n9049);
   U5799 : OAI22_X1 port map( A1 => n20486, A2 => n20278, B1 => n3459, B2 => 
                           n20284, ZN => n9050);
   U5800 : OAI22_X1 port map( A1 => n20489, A2 => n20277, B1 => n3458, B2 => 
                           n20283, ZN => n9051);
   U5801 : OAI22_X1 port map( A1 => n20492, A2 => n20276, B1 => n3457, B2 => 
                           n20283, ZN => n9052);
   U5802 : OAI22_X1 port map( A1 => n20495, A2 => n20278, B1 => n3456, B2 => 
                           n20283, ZN => n9053);
   U5803 : OAI22_X1 port map( A1 => n20498, A2 => n20277, B1 => n3455, B2 => 
                           n20283, ZN => n9054);
   U5804 : OAI22_X1 port map( A1 => n20501, A2 => n20276, B1 => n3454, B2 => 
                           n20282, ZN => n9055);
   U5805 : OAI22_X1 port map( A1 => n20504, A2 => n20278, B1 => n3453, B2 => 
                           n20282, ZN => n9056);
   U5806 : OAI22_X1 port map( A1 => n20507, A2 => n20277, B1 => n3452, B2 => 
                           n20282, ZN => n9057);
   U5807 : OAI22_X1 port map( A1 => n20510, A2 => n20277, B1 => n3451, B2 => 
                           n20282, ZN => n9058);
   U5808 : OAI22_X1 port map( A1 => n20513, A2 => n20278, B1 => n3450, B2 => 
                           n20281, ZN => n9059);
   U5809 : OAI22_X1 port map( A1 => n20516, A2 => n20277, B1 => n3449, B2 => 
                           n20281, ZN => n9060);
   U5810 : OAI22_X1 port map( A1 => n20519, A2 => n20276, B1 => n3448, B2 => 
                           n20281, ZN => n9061);
   U5811 : OAI22_X1 port map( A1 => n20522, A2 => n20276, B1 => n3447, B2 => 
                           n20281, ZN => n9062);
   U5812 : OAI22_X1 port map( A1 => n20525, A2 => n20278, B1 => n3446, B2 => 
                           n20280, ZN => n9063);
   U5813 : OAI22_X1 port map( A1 => n20528, A2 => n20277, B1 => n3445, B2 => 
                           n20280, ZN => n9064);
   U5814 : OAI22_X1 port map( A1 => n20531, A2 => n20276, B1 => n3444, B2 => 
                           n20280, ZN => n9065);
   U5815 : OAI22_X1 port map( A1 => n20534, A2 => n20278, B1 => n3443, B2 => 
                           n20280, ZN => n9066);
   U5816 : OAI22_X1 port map( A1 => n20537, A2 => n20278, B1 => n3442, B2 => 
                           n20279, ZN => n9067);
   U5817 : OAI22_X1 port map( A1 => n20540, A2 => n20277, B1 => n3441, B2 => 
                           n20279, ZN => n9068);
   U5818 : OAI22_X1 port map( A1 => n20543, A2 => n20276, B1 => n3440, B2 => 
                           n20279, ZN => n9069);
   U5819 : OAI22_X1 port map( A1 => n20574, A2 => n20277, B1 => n3439, B2 => 
                           n20279, ZN => n9070);
   U5820 : OAI22_X1 port map( A1 => n20357, A2 => n20277, B1 => n3502, B2 => 
                           n20294, ZN => n9007);
   U5821 : OAI22_X1 port map( A1 => n20360, A2 => n20276, B1 => n3501, B2 => 
                           n20294, ZN => n9008);
   U5822 : OAI22_X1 port map( A1 => n20363, A2 => n20276, B1 => n3500, B2 => 
                           n20294, ZN => n9009);
   U5823 : OAI22_X1 port map( A1 => n20366, A2 => n20278, B1 => n3499, B2 => 
                           n20294, ZN => n9010);
   U5824 : OAI22_X1 port map( A1 => n20391, A2 => n19634, B1 => n5041, B2 => 
                           n19647, ZN => n7547);
   U5825 : OAI22_X1 port map( A1 => n20394, A2 => n19633, B1 => n5040, B2 => 
                           n19647, ZN => n7548);
   U5826 : OAI22_X1 port map( A1 => n20397, A2 => n19632, B1 => n5039, B2 => 
                           n19647, ZN => n7549);
   U5827 : OAI22_X1 port map( A1 => n20400, A2 => n19634, B1 => n5038, B2 => 
                           n19647, ZN => n7550);
   U5828 : OAI22_X1 port map( A1 => n20403, A2 => n19634, B1 => n5037, B2 => 
                           n19646, ZN => n7551);
   U5829 : OAI22_X1 port map( A1 => n20406, A2 => n19634, B1 => n5036, B2 => 
                           n19646, ZN => n7552);
   U5830 : OAI22_X1 port map( A1 => n20409, A2 => n19634, B1 => n5035, B2 => 
                           n19646, ZN => n7553);
   U5831 : OAI22_X1 port map( A1 => n20412, A2 => n19634, B1 => n5034, B2 => 
                           n19646, ZN => n7554);
   U5832 : OAI22_X1 port map( A1 => n20415, A2 => n19634, B1 => n5033, B2 => 
                           n19645, ZN => n7555);
   U5833 : OAI22_X1 port map( A1 => n20418, A2 => n19634, B1 => n5032, B2 => 
                           n19645, ZN => n7556);
   U5834 : OAI22_X1 port map( A1 => n20421, A2 => n19634, B1 => n5031, B2 => 
                           n19645, ZN => n7557);
   U5835 : OAI22_X1 port map( A1 => n20424, A2 => n19634, B1 => n5030, B2 => 
                           n19645, ZN => n7558);
   U5836 : OAI22_X1 port map( A1 => n20427, A2 => n19634, B1 => n5029, B2 => 
                           n19644, ZN => n7559);
   U5837 : OAI22_X1 port map( A1 => n20430, A2 => n19634, B1 => n5028, B2 => 
                           n19644, ZN => n7560);
   U5838 : OAI22_X1 port map( A1 => n20433, A2 => n19634, B1 => n5027, B2 => 
                           n19644, ZN => n7561);
   U5839 : OAI22_X1 port map( A1 => n20436, A2 => n19634, B1 => n5026, B2 => 
                           n19644, ZN => n7562);
   U5840 : OAI22_X1 port map( A1 => n20439, A2 => n19633, B1 => n5025, B2 => 
                           n19643, ZN => n7563);
   U5841 : OAI22_X1 port map( A1 => n20442, A2 => n19633, B1 => n5024, B2 => 
                           n19643, ZN => n7564);
   U5842 : OAI22_X1 port map( A1 => n20445, A2 => n19633, B1 => n5023, B2 => 
                           n19643, ZN => n7565);
   U5843 : OAI22_X1 port map( A1 => n20448, A2 => n19633, B1 => n5022, B2 => 
                           n19643, ZN => n7566);
   U5844 : OAI22_X1 port map( A1 => n20451, A2 => n19633, B1 => n5021, B2 => 
                           n19642, ZN => n7567);
   U5845 : OAI22_X1 port map( A1 => n20454, A2 => n19633, B1 => n5020, B2 => 
                           n19642, ZN => n7568);
   U5846 : OAI22_X1 port map( A1 => n20457, A2 => n19633, B1 => n5019, B2 => 
                           n19642, ZN => n7569);
   U5847 : OAI22_X1 port map( A1 => n20460, A2 => n19633, B1 => n5018, B2 => 
                           n19642, ZN => n7570);
   U5848 : OAI22_X1 port map( A1 => n20463, A2 => n19633, B1 => n5017, B2 => 
                           n19641, ZN => n7571);
   U5849 : OAI22_X1 port map( A1 => n20466, A2 => n19633, B1 => n5016, B2 => 
                           n19641, ZN => n7572);
   U5850 : OAI22_X1 port map( A1 => n20469, A2 => n19633, B1 => n5015, B2 => 
                           n19641, ZN => n7573);
   U5851 : OAI22_X1 port map( A1 => n20472, A2 => n19633, B1 => n5014, B2 => 
                           n19641, ZN => n7574);
   U5852 : OAI22_X1 port map( A1 => n20475, A2 => n19632, B1 => n5013, B2 => 
                           n19640, ZN => n7575);
   U5853 : OAI22_X1 port map( A1 => n20478, A2 => n19632, B1 => n5012, B2 => 
                           n19640, ZN => n7576);
   U5854 : OAI22_X1 port map( A1 => n20481, A2 => n19632, B1 => n5011, B2 => 
                           n19640, ZN => n7577);
   U5855 : OAI22_X1 port map( A1 => n20484, A2 => n19632, B1 => n5010, B2 => 
                           n19640, ZN => n7578);
   U5856 : OAI22_X1 port map( A1 => n20487, A2 => n19632, B1 => n5009, B2 => 
                           n19639, ZN => n7579);
   U5857 : OAI22_X1 port map( A1 => n20490, A2 => n19632, B1 => n5008, B2 => 
                           n19639, ZN => n7580);
   U5858 : OAI22_X1 port map( A1 => n20493, A2 => n19632, B1 => n5007, B2 => 
                           n19639, ZN => n7581);
   U5859 : OAI22_X1 port map( A1 => n20496, A2 => n19632, B1 => n5006, B2 => 
                           n19639, ZN => n7582);
   U5860 : OAI22_X1 port map( A1 => n20499, A2 => n19632, B1 => n5005, B2 => 
                           n19638, ZN => n7583);
   U5861 : OAI22_X1 port map( A1 => n20502, A2 => n19632, B1 => n5004, B2 => 
                           n19638, ZN => n7584);
   U5862 : OAI22_X1 port map( A1 => n20505, A2 => n19632, B1 => n5003, B2 => 
                           n19638, ZN => n7585);
   U5863 : OAI22_X1 port map( A1 => n20508, A2 => n19632, B1 => n5002, B2 => 
                           n19638, ZN => n7586);
   U5864 : OAI22_X1 port map( A1 => n20511, A2 => n19632, B1 => n5001, B2 => 
                           n19637, ZN => n7587);
   U5865 : OAI22_X1 port map( A1 => n20514, A2 => n19634, B1 => n5000, B2 => 
                           n19637, ZN => n7588);
   U5866 : OAI22_X1 port map( A1 => n20517, A2 => n19633, B1 => n4999, B2 => 
                           n19637, ZN => n7589);
   U5867 : OAI22_X1 port map( A1 => n20520, A2 => n19632, B1 => n4998, B2 => 
                           n19637, ZN => n7590);
   U5868 : OAI22_X1 port map( A1 => n20523, A2 => n19634, B1 => n4997, B2 => 
                           n19636, ZN => n7591);
   U5869 : OAI22_X1 port map( A1 => n20526, A2 => n19634, B1 => n4996, B2 => 
                           n19636, ZN => n7592);
   U5870 : OAI22_X1 port map( A1 => n20529, A2 => n19633, B1 => n4995, B2 => 
                           n19636, ZN => n7593);
   U5871 : OAI22_X1 port map( A1 => n20532, A2 => n19632, B1 => n4994, B2 => 
                           n19636, ZN => n7594);
   U5872 : OAI22_X1 port map( A1 => n20535, A2 => n19633, B1 => n4993, B2 => 
                           n19635, ZN => n7595);
   U5873 : OAI22_X1 port map( A1 => n20538, A2 => n19634, B1 => n4992, B2 => 
                           n19635, ZN => n7596);
   U5874 : OAI22_X1 port map( A1 => n20541, A2 => n19633, B1 => n4991, B2 => 
                           n19635, ZN => n7597);
   U5875 : OAI22_X1 port map( A1 => n20572, A2 => n19632, B1 => n4990, B2 => 
                           n19635, ZN => n7598);
   U5876 : OAI22_X1 port map( A1 => n20367, A2 => n19746, B1 => n4779, B2 => 
                           n19761, ZN => n7795);
   U5877 : OAI22_X1 port map( A1 => n20370, A2 => n19746, B1 => n4778, B2 => 
                           n19761, ZN => n7796);
   U5878 : OAI22_X1 port map( A1 => n20373, A2 => n19746, B1 => n4777, B2 => 
                           n19761, ZN => n7797);
   U5879 : OAI22_X1 port map( A1 => n20376, A2 => n19746, B1 => n4776, B2 => 
                           n19761, ZN => n7798);
   U5880 : OAI22_X1 port map( A1 => n20379, A2 => n19746, B1 => n4775, B2 => 
                           n19760, ZN => n7799);
   U5881 : OAI22_X1 port map( A1 => n20382, A2 => n19746, B1 => n4774, B2 => 
                           n19760, ZN => n7800);
   U5882 : OAI22_X1 port map( A1 => n20385, A2 => n19746, B1 => n4773, B2 => 
                           n19760, ZN => n7801);
   U5883 : OAI22_X1 port map( A1 => n20388, A2 => n19746, B1 => n4772, B2 => 
                           n19760, ZN => n7802);
   U5884 : OAI22_X1 port map( A1 => n20391, A2 => n19746, B1 => n4771, B2 => 
                           n19759, ZN => n7803);
   U5885 : OAI22_X1 port map( A1 => n20394, A2 => n19746, B1 => n4770, B2 => 
                           n19759, ZN => n7804);
   U5886 : OAI22_X1 port map( A1 => n20397, A2 => n19746, B1 => n4769, B2 => 
                           n19759, ZN => n7805);
   U5887 : OAI22_X1 port map( A1 => n20400, A2 => n19746, B1 => n4768, B2 => 
                           n19759, ZN => n7806);
   U5888 : OAI22_X1 port map( A1 => n20403, A2 => n19745, B1 => n4767, B2 => 
                           n19758, ZN => n7807);
   U5889 : OAI22_X1 port map( A1 => n20406, A2 => n19745, B1 => n4766, B2 => 
                           n19758, ZN => n7808);
   U5890 : OAI22_X1 port map( A1 => n20409, A2 => n19745, B1 => n4765, B2 => 
                           n19758, ZN => n7809);
   U5891 : OAI22_X1 port map( A1 => n20412, A2 => n19745, B1 => n4764, B2 => 
                           n19758, ZN => n7810);
   U5892 : OAI22_X1 port map( A1 => n20415, A2 => n19745, B1 => n4763, B2 => 
                           n19757, ZN => n7811);
   U5893 : OAI22_X1 port map( A1 => n20418, A2 => n19745, B1 => n4762, B2 => 
                           n19757, ZN => n7812);
   U5894 : OAI22_X1 port map( A1 => n20421, A2 => n19745, B1 => n4761, B2 => 
                           n19757, ZN => n7813);
   U5895 : OAI22_X1 port map( A1 => n20424, A2 => n19745, B1 => n4760, B2 => 
                           n19757, ZN => n7814);
   U5896 : OAI22_X1 port map( A1 => n20427, A2 => n19745, B1 => n4759, B2 => 
                           n19756, ZN => n7815);
   U5897 : OAI22_X1 port map( A1 => n20430, A2 => n19745, B1 => n4758, B2 => 
                           n19756, ZN => n7816);
   U5898 : OAI22_X1 port map( A1 => n20433, A2 => n19745, B1 => n4757, B2 => 
                           n19756, ZN => n7817);
   U5899 : OAI22_X1 port map( A1 => n20436, A2 => n19745, B1 => n4756, B2 => 
                           n19756, ZN => n7818);
   U5900 : OAI22_X1 port map( A1 => n20439, A2 => n19744, B1 => n4755, B2 => 
                           n19755, ZN => n7819);
   U5901 : OAI22_X1 port map( A1 => n20442, A2 => n19744, B1 => n4754, B2 => 
                           n19755, ZN => n7820);
   U5902 : OAI22_X1 port map( A1 => n20445, A2 => n19744, B1 => n4753, B2 => 
                           n19755, ZN => n7821);
   U5903 : OAI22_X1 port map( A1 => n20448, A2 => n19744, B1 => n4752, B2 => 
                           n19755, ZN => n7822);
   U5904 : OAI22_X1 port map( A1 => n20451, A2 => n19744, B1 => n4751, B2 => 
                           n19754, ZN => n7823);
   U5905 : OAI22_X1 port map( A1 => n20454, A2 => n19744, B1 => n4750, B2 => 
                           n19754, ZN => n7824);
   U5906 : OAI22_X1 port map( A1 => n20457, A2 => n19744, B1 => n4749, B2 => 
                           n19754, ZN => n7825);
   U5907 : OAI22_X1 port map( A1 => n20460, A2 => n19744, B1 => n4748, B2 => 
                           n19754, ZN => n7826);
   U5908 : OAI22_X1 port map( A1 => n20463, A2 => n19744, B1 => n4747, B2 => 
                           n19753, ZN => n7827);
   U5909 : OAI22_X1 port map( A1 => n20466, A2 => n19744, B1 => n4746, B2 => 
                           n19753, ZN => n7828);
   U5910 : OAI22_X1 port map( A1 => n20469, A2 => n19744, B1 => n4745, B2 => 
                           n19753, ZN => n7829);
   U5911 : OAI22_X1 port map( A1 => n20472, A2 => n19744, B1 => n4744, B2 => 
                           n19753, ZN => n7830);
   U5912 : OAI22_X1 port map( A1 => n20475, A2 => n19746, B1 => n4743, B2 => 
                           n19752, ZN => n7831);
   U5913 : OAI22_X1 port map( A1 => n20478, A2 => n19745, B1 => n4742, B2 => 
                           n19752, ZN => n7832);
   U5914 : OAI22_X1 port map( A1 => n20481, A2 => n19744, B1 => n4741, B2 => 
                           n19752, ZN => n7833);
   U5915 : OAI22_X1 port map( A1 => n20484, A2 => n19746, B1 => n4740, B2 => 
                           n19752, ZN => n7834);
   U5916 : OAI22_X1 port map( A1 => n20487, A2 => n19745, B1 => n4739, B2 => 
                           n19751, ZN => n7835);
   U5917 : OAI22_X1 port map( A1 => n20490, A2 => n19744, B1 => n4738, B2 => 
                           n19751, ZN => n7836);
   U5918 : OAI22_X1 port map( A1 => n20493, A2 => n19746, B1 => n4737, B2 => 
                           n19751, ZN => n7837);
   U5919 : OAI22_X1 port map( A1 => n20496, A2 => n19745, B1 => n4736, B2 => 
                           n19751, ZN => n7838);
   U5920 : OAI22_X1 port map( A1 => n20499, A2 => n19744, B1 => n4735, B2 => 
                           n19750, ZN => n7839);
   U5921 : OAI22_X1 port map( A1 => n20502, A2 => n19746, B1 => n4734, B2 => 
                           n19750, ZN => n7840);
   U5922 : OAI22_X1 port map( A1 => n20505, A2 => n19745, B1 => n4733, B2 => 
                           n19750, ZN => n7841);
   U5923 : OAI22_X1 port map( A1 => n20508, A2 => n19745, B1 => n4732, B2 => 
                           n19750, ZN => n7842);
   U5924 : OAI22_X1 port map( A1 => n20511, A2 => n19746, B1 => n4731, B2 => 
                           n19749, ZN => n7843);
   U5925 : OAI22_X1 port map( A1 => n20514, A2 => n19745, B1 => n4730, B2 => 
                           n19749, ZN => n7844);
   U5926 : OAI22_X1 port map( A1 => n20517, A2 => n19744, B1 => n4729, B2 => 
                           n19749, ZN => n7845);
   U5927 : OAI22_X1 port map( A1 => n20520, A2 => n19744, B1 => n4728, B2 => 
                           n19749, ZN => n7846);
   U5928 : OAI22_X1 port map( A1 => n20523, A2 => n19746, B1 => n4727, B2 => 
                           n19748, ZN => n7847);
   U5929 : OAI22_X1 port map( A1 => n20526, A2 => n19745, B1 => n4726, B2 => 
                           n19748, ZN => n7848);
   U5930 : OAI22_X1 port map( A1 => n20529, A2 => n19744, B1 => n4725, B2 => 
                           n19748, ZN => n7849);
   U5931 : OAI22_X1 port map( A1 => n20532, A2 => n19746, B1 => n4724, B2 => 
                           n19748, ZN => n7850);
   U5932 : OAI22_X1 port map( A1 => n20535, A2 => n19746, B1 => n4723, B2 => 
                           n19747, ZN => n7851);
   U5933 : OAI22_X1 port map( A1 => n20538, A2 => n19745, B1 => n4722, B2 => 
                           n19747, ZN => n7852);
   U5934 : OAI22_X1 port map( A1 => n20541, A2 => n19744, B1 => n4721, B2 => 
                           n19747, ZN => n7853);
   U5935 : OAI22_X1 port map( A1 => n20572, A2 => n19745, B1 => n4720, B2 => 
                           n19747, ZN => n7854);
   U5936 : OAI22_X1 port map( A1 => n20355, A2 => n19745, B1 => n4783, B2 => 
                           n19762, ZN => n7791);
   U5937 : OAI22_X1 port map( A1 => n20358, A2 => n19744, B1 => n4782, B2 => 
                           n19762, ZN => n7792);
   U5938 : OAI22_X1 port map( A1 => n20361, A2 => n19744, B1 => n4781, B2 => 
                           n19762, ZN => n7793);
   U5939 : OAI22_X1 port map( A1 => n20364, A2 => n19746, B1 => n4780, B2 => 
                           n19762, ZN => n7794);
   U5940 : OAI22_X1 port map( A1 => n20391, A2 => n19662, B1 => n4975, B2 => 
                           n19675, ZN => n7611);
   U5941 : OAI22_X1 port map( A1 => n20394, A2 => n19661, B1 => n4974, B2 => 
                           n19675, ZN => n7612);
   U5942 : OAI22_X1 port map( A1 => n20397, A2 => n19660, B1 => n4973, B2 => 
                           n19675, ZN => n7613);
   U5943 : OAI22_X1 port map( A1 => n20400, A2 => n19662, B1 => n4972, B2 => 
                           n19675, ZN => n7614);
   U5944 : OAI22_X1 port map( A1 => n20403, A2 => n19662, B1 => n4971, B2 => 
                           n19674, ZN => n7615);
   U5945 : OAI22_X1 port map( A1 => n20406, A2 => n19662, B1 => n4970, B2 => 
                           n19674, ZN => n7616);
   U5946 : OAI22_X1 port map( A1 => n20409, A2 => n19662, B1 => n4969, B2 => 
                           n19674, ZN => n7617);
   U5947 : OAI22_X1 port map( A1 => n20412, A2 => n19662, B1 => n4968, B2 => 
                           n19674, ZN => n7618);
   U5948 : OAI22_X1 port map( A1 => n20415, A2 => n19662, B1 => n4967, B2 => 
                           n19673, ZN => n7619);
   U5949 : OAI22_X1 port map( A1 => n20418, A2 => n19662, B1 => n4966, B2 => 
                           n19673, ZN => n7620);
   U5950 : OAI22_X1 port map( A1 => n20421, A2 => n19662, B1 => n4965, B2 => 
                           n19673, ZN => n7621);
   U5951 : OAI22_X1 port map( A1 => n20424, A2 => n19662, B1 => n4964, B2 => 
                           n19673, ZN => n7622);
   U5952 : OAI22_X1 port map( A1 => n20427, A2 => n19662, B1 => n4963, B2 => 
                           n19672, ZN => n7623);
   U5953 : OAI22_X1 port map( A1 => n20430, A2 => n19662, B1 => n4962, B2 => 
                           n19672, ZN => n7624);
   U5954 : OAI22_X1 port map( A1 => n20433, A2 => n19662, B1 => n4961, B2 => 
                           n19672, ZN => n7625);
   U5955 : OAI22_X1 port map( A1 => n20436, A2 => n19662, B1 => n4960, B2 => 
                           n19672, ZN => n7626);
   U5956 : OAI22_X1 port map( A1 => n20439, A2 => n19661, B1 => n4959, B2 => 
                           n19671, ZN => n7627);
   U5957 : OAI22_X1 port map( A1 => n20442, A2 => n19661, B1 => n4958, B2 => 
                           n19671, ZN => n7628);
   U5958 : OAI22_X1 port map( A1 => n20445, A2 => n19661, B1 => n4957, B2 => 
                           n19671, ZN => n7629);
   U5959 : OAI22_X1 port map( A1 => n20448, A2 => n19661, B1 => n4956, B2 => 
                           n19671, ZN => n7630);
   U5960 : OAI22_X1 port map( A1 => n20451, A2 => n19661, B1 => n4955, B2 => 
                           n19670, ZN => n7631);
   U5961 : OAI22_X1 port map( A1 => n20454, A2 => n19661, B1 => n4954, B2 => 
                           n19670, ZN => n7632);
   U5962 : OAI22_X1 port map( A1 => n20457, A2 => n19661, B1 => n4953, B2 => 
                           n19670, ZN => n7633);
   U5963 : OAI22_X1 port map( A1 => n20460, A2 => n19661, B1 => n4952, B2 => 
                           n19670, ZN => n7634);
   U5964 : OAI22_X1 port map( A1 => n20463, A2 => n19661, B1 => n4951, B2 => 
                           n19669, ZN => n7635);
   U5965 : OAI22_X1 port map( A1 => n20466, A2 => n19661, B1 => n4950, B2 => 
                           n19669, ZN => n7636);
   U5966 : OAI22_X1 port map( A1 => n20469, A2 => n19661, B1 => n4949, B2 => 
                           n19669, ZN => n7637);
   U5967 : OAI22_X1 port map( A1 => n20472, A2 => n19661, B1 => n4948, B2 => 
                           n19669, ZN => n7638);
   U5968 : OAI22_X1 port map( A1 => n20475, A2 => n19660, B1 => n4947, B2 => 
                           n19668, ZN => n7639);
   U5969 : OAI22_X1 port map( A1 => n20478, A2 => n19660, B1 => n4946, B2 => 
                           n19668, ZN => n7640);
   U5970 : OAI22_X1 port map( A1 => n20481, A2 => n19660, B1 => n4945, B2 => 
                           n19668, ZN => n7641);
   U5971 : OAI22_X1 port map( A1 => n20484, A2 => n19660, B1 => n4944, B2 => 
                           n19668, ZN => n7642);
   U5972 : OAI22_X1 port map( A1 => n20487, A2 => n19660, B1 => n4943, B2 => 
                           n19667, ZN => n7643);
   U5973 : OAI22_X1 port map( A1 => n20490, A2 => n19660, B1 => n4942, B2 => 
                           n19667, ZN => n7644);
   U5974 : OAI22_X1 port map( A1 => n20493, A2 => n19660, B1 => n4941, B2 => 
                           n19667, ZN => n7645);
   U5975 : OAI22_X1 port map( A1 => n20496, A2 => n19660, B1 => n4940, B2 => 
                           n19667, ZN => n7646);
   U5976 : OAI22_X1 port map( A1 => n20499, A2 => n19660, B1 => n4939, B2 => 
                           n19666, ZN => n7647);
   U5977 : OAI22_X1 port map( A1 => n20502, A2 => n19660, B1 => n4938, B2 => 
                           n19666, ZN => n7648);
   U5978 : OAI22_X1 port map( A1 => n20505, A2 => n19660, B1 => n4937, B2 => 
                           n19666, ZN => n7649);
   U5979 : OAI22_X1 port map( A1 => n20508, A2 => n19660, B1 => n4936, B2 => 
                           n19666, ZN => n7650);
   U5980 : OAI22_X1 port map( A1 => n20511, A2 => n19660, B1 => n4935, B2 => 
                           n19665, ZN => n7651);
   U5981 : OAI22_X1 port map( A1 => n20514, A2 => n19662, B1 => n4934, B2 => 
                           n19665, ZN => n7652);
   U5982 : OAI22_X1 port map( A1 => n20517, A2 => n19661, B1 => n4933, B2 => 
                           n19665, ZN => n7653);
   U5983 : OAI22_X1 port map( A1 => n20520, A2 => n19660, B1 => n4932, B2 => 
                           n19665, ZN => n7654);
   U5984 : OAI22_X1 port map( A1 => n20523, A2 => n19662, B1 => n4931, B2 => 
                           n19664, ZN => n7655);
   U5985 : OAI22_X1 port map( A1 => n20526, A2 => n19662, B1 => n4930, B2 => 
                           n19664, ZN => n7656);
   U5986 : OAI22_X1 port map( A1 => n20529, A2 => n19661, B1 => n4929, B2 => 
                           n19664, ZN => n7657);
   U5987 : OAI22_X1 port map( A1 => n20532, A2 => n19660, B1 => n4928, B2 => 
                           n19664, ZN => n7658);
   U5988 : OAI22_X1 port map( A1 => n20535, A2 => n19661, B1 => n4927, B2 => 
                           n19663, ZN => n7659);
   U5989 : OAI22_X1 port map( A1 => n20538, A2 => n19662, B1 => n4926, B2 => 
                           n19663, ZN => n7660);
   U5990 : OAI22_X1 port map( A1 => n20541, A2 => n19661, B1 => n4925, B2 => 
                           n19663, ZN => n7661);
   U5991 : OAI22_X1 port map( A1 => n20572, A2 => n19660, B1 => n4924, B2 => 
                           n19663, ZN => n7662);
   U5992 : OAI22_X1 port map( A1 => n20367, A2 => n19661, B1 => n4983, B2 => 
                           n19677, ZN => n7603);
   U5993 : OAI22_X1 port map( A1 => n20370, A2 => n19660, B1 => n4982, B2 => 
                           n19677, ZN => n7604);
   U5994 : OAI22_X1 port map( A1 => n20373, A2 => n19662, B1 => n4981, B2 => 
                           n19677, ZN => n7605);
   U5995 : OAI22_X1 port map( A1 => n20376, A2 => n19661, B1 => n4980, B2 => 
                           n19677, ZN => n7606);
   U5996 : OAI22_X1 port map( A1 => n20379, A2 => n19660, B1 => n4979, B2 => 
                           n19676, ZN => n7607);
   U5997 : OAI22_X1 port map( A1 => n20382, A2 => n19662, B1 => n4978, B2 => 
                           n19676, ZN => n7608);
   U5998 : OAI22_X1 port map( A1 => n20385, A2 => n19661, B1 => n4977, B2 => 
                           n19676, ZN => n7609);
   U5999 : OAI22_X1 port map( A1 => n20388, A2 => n19661, B1 => n4976, B2 => 
                           n19676, ZN => n7610);
   U6000 : OAI22_X1 port map( A1 => n20355, A2 => n19662, B1 => n4987, B2 => 
                           n19678, ZN => n7599);
   U6001 : OAI22_X1 port map( A1 => n20358, A2 => n19661, B1 => n4986, B2 => 
                           n19678, ZN => n7600);
   U6002 : OAI22_X1 port map( A1 => n20361, A2 => n19660, B1 => n4985, B2 => 
                           n19678, ZN => n7601);
   U6003 : OAI22_X1 port map( A1 => n20364, A2 => n19660, B1 => n4984, B2 => 
                           n19678, ZN => n7602);
   U6004 : OAI22_X1 port map( A1 => n20367, A2 => n19633, B1 => n5049, B2 => 
                           n19649, ZN => n7539);
   U6005 : OAI22_X1 port map( A1 => n20370, A2 => n19632, B1 => n5048, B2 => 
                           n19649, ZN => n7540);
   U6006 : OAI22_X1 port map( A1 => n20373, A2 => n19634, B1 => n5047, B2 => 
                           n19649, ZN => n7541);
   U6007 : OAI22_X1 port map( A1 => n20376, A2 => n19633, B1 => n5046, B2 => 
                           n19649, ZN => n7542);
   U6008 : OAI22_X1 port map( A1 => n20379, A2 => n19632, B1 => n5045, B2 => 
                           n19648, ZN => n7543);
   U6009 : OAI22_X1 port map( A1 => n20382, A2 => n19634, B1 => n5044, B2 => 
                           n19648, ZN => n7544);
   U6010 : OAI22_X1 port map( A1 => n20385, A2 => n19633, B1 => n5043, B2 => 
                           n19648, ZN => n7545);
   U6011 : OAI22_X1 port map( A1 => n20388, A2 => n19633, B1 => n5042, B2 => 
                           n19648, ZN => n7546);
   U6012 : OAI22_X1 port map( A1 => n20355, A2 => n19634, B1 => n5053, B2 => 
                           n19650, ZN => n7535);
   U6013 : OAI22_X1 port map( A1 => n20358, A2 => n19633, B1 => n5052, B2 => 
                           n19650, ZN => n7536);
   U6014 : OAI22_X1 port map( A1 => n20361, A2 => n19632, B1 => n5051, B2 => 
                           n19650, ZN => n7537);
   U6015 : OAI22_X1 port map( A1 => n20364, A2 => n19632, B1 => n5050, B2 => 
                           n19650, ZN => n7538);
   U6016 : OAI22_X1 port map( A1 => n20368, A2 => n20054, B1 => n4033, B2 => 
                           n20069, ZN => n8499);
   U6017 : OAI22_X1 port map( A1 => n20371, A2 => n20054, B1 => n4032, B2 => 
                           n20069, ZN => n8500);
   U6018 : OAI22_X1 port map( A1 => n20374, A2 => n20054, B1 => n4031, B2 => 
                           n20069, ZN => n8501);
   U6019 : OAI22_X1 port map( A1 => n20377, A2 => n20054, B1 => n4030, B2 => 
                           n20069, ZN => n8502);
   U6020 : OAI22_X1 port map( A1 => n20380, A2 => n20054, B1 => n4029, B2 => 
                           n20068, ZN => n8503);
   U6021 : OAI22_X1 port map( A1 => n20383, A2 => n20054, B1 => n4028, B2 => 
                           n20068, ZN => n8504);
   U6022 : OAI22_X1 port map( A1 => n20386, A2 => n20054, B1 => n4027, B2 => 
                           n20068, ZN => n8505);
   U6023 : OAI22_X1 port map( A1 => n20389, A2 => n20054, B1 => n4026, B2 => 
                           n20068, ZN => n8506);
   U6024 : OAI22_X1 port map( A1 => n20392, A2 => n20054, B1 => n4025, B2 => 
                           n20067, ZN => n8507);
   U6025 : OAI22_X1 port map( A1 => n20395, A2 => n20054, B1 => n4024, B2 => 
                           n20067, ZN => n8508);
   U6026 : OAI22_X1 port map( A1 => n20398, A2 => n20054, B1 => n4023, B2 => 
                           n20067, ZN => n8509);
   U6027 : OAI22_X1 port map( A1 => n20401, A2 => n20054, B1 => n4022, B2 => 
                           n20067, ZN => n8510);
   U6028 : OAI22_X1 port map( A1 => n20404, A2 => n20053, B1 => n4021, B2 => 
                           n20066, ZN => n8511);
   U6029 : OAI22_X1 port map( A1 => n20407, A2 => n20053, B1 => n4020, B2 => 
                           n20066, ZN => n8512);
   U6030 : OAI22_X1 port map( A1 => n20410, A2 => n20053, B1 => n4019, B2 => 
                           n20066, ZN => n8513);
   U6031 : OAI22_X1 port map( A1 => n20413, A2 => n20053, B1 => n4018, B2 => 
                           n20066, ZN => n8514);
   U6032 : OAI22_X1 port map( A1 => n20416, A2 => n20053, B1 => n4017, B2 => 
                           n20065, ZN => n8515);
   U6033 : OAI22_X1 port map( A1 => n20419, A2 => n20053, B1 => n4016, B2 => 
                           n20065, ZN => n8516);
   U6034 : OAI22_X1 port map( A1 => n20422, A2 => n20053, B1 => n4015, B2 => 
                           n20065, ZN => n8517);
   U6035 : OAI22_X1 port map( A1 => n20425, A2 => n20053, B1 => n4014, B2 => 
                           n20065, ZN => n8518);
   U6036 : OAI22_X1 port map( A1 => n20428, A2 => n20053, B1 => n4013, B2 => 
                           n20064, ZN => n8519);
   U6037 : OAI22_X1 port map( A1 => n20431, A2 => n20053, B1 => n4012, B2 => 
                           n20064, ZN => n8520);
   U6038 : OAI22_X1 port map( A1 => n20434, A2 => n20053, B1 => n4011, B2 => 
                           n20064, ZN => n8521);
   U6039 : OAI22_X1 port map( A1 => n20437, A2 => n20053, B1 => n4010, B2 => 
                           n20064, ZN => n8522);
   U6040 : OAI22_X1 port map( A1 => n20440, A2 => n20052, B1 => n4009, B2 => 
                           n20063, ZN => n8523);
   U6041 : OAI22_X1 port map( A1 => n20443, A2 => n20052, B1 => n4008, B2 => 
                           n20063, ZN => n8524);
   U6042 : OAI22_X1 port map( A1 => n20446, A2 => n20052, B1 => n4007, B2 => 
                           n20063, ZN => n8525);
   U6043 : OAI22_X1 port map( A1 => n20449, A2 => n20052, B1 => n4006, B2 => 
                           n20063, ZN => n8526);
   U6044 : OAI22_X1 port map( A1 => n20452, A2 => n20052, B1 => n4005, B2 => 
                           n20062, ZN => n8527);
   U6045 : OAI22_X1 port map( A1 => n20455, A2 => n20052, B1 => n4004, B2 => 
                           n20062, ZN => n8528);
   U6046 : OAI22_X1 port map( A1 => n20458, A2 => n20052, B1 => n4003, B2 => 
                           n20062, ZN => n8529);
   U6047 : OAI22_X1 port map( A1 => n20461, A2 => n20052, B1 => n4002, B2 => 
                           n20062, ZN => n8530);
   U6048 : OAI22_X1 port map( A1 => n20464, A2 => n20052, B1 => n4001, B2 => 
                           n20061, ZN => n8531);
   U6049 : OAI22_X1 port map( A1 => n20467, A2 => n20052, B1 => n4000, B2 => 
                           n20061, ZN => n8532);
   U6050 : OAI22_X1 port map( A1 => n20470, A2 => n20052, B1 => n3999, B2 => 
                           n20061, ZN => n8533);
   U6051 : OAI22_X1 port map( A1 => n20473, A2 => n20052, B1 => n3998, B2 => 
                           n20061, ZN => n8534);
   U6052 : OAI22_X1 port map( A1 => n20476, A2 => n20054, B1 => n3997, B2 => 
                           n20060, ZN => n8535);
   U6053 : OAI22_X1 port map( A1 => n20479, A2 => n20053, B1 => n3996, B2 => 
                           n20060, ZN => n8536);
   U6054 : OAI22_X1 port map( A1 => n20482, A2 => n20052, B1 => n3995, B2 => 
                           n20060, ZN => n8537);
   U6055 : OAI22_X1 port map( A1 => n20485, A2 => n20054, B1 => n3994, B2 => 
                           n20060, ZN => n8538);
   U6056 : OAI22_X1 port map( A1 => n20488, A2 => n20053, B1 => n3993, B2 => 
                           n20059, ZN => n8539);
   U6057 : OAI22_X1 port map( A1 => n20491, A2 => n20052, B1 => n3992, B2 => 
                           n20059, ZN => n8540);
   U6058 : OAI22_X1 port map( A1 => n20494, A2 => n20054, B1 => n3991, B2 => 
                           n20059, ZN => n8541);
   U6059 : OAI22_X1 port map( A1 => n20497, A2 => n20053, B1 => n3990, B2 => 
                           n20059, ZN => n8542);
   U6060 : OAI22_X1 port map( A1 => n20500, A2 => n20052, B1 => n3989, B2 => 
                           n20058, ZN => n8543);
   U6061 : OAI22_X1 port map( A1 => n20503, A2 => n20054, B1 => n3988, B2 => 
                           n20058, ZN => n8544);
   U6062 : OAI22_X1 port map( A1 => n20506, A2 => n20053, B1 => n3987, B2 => 
                           n20058, ZN => n8545);
   U6063 : OAI22_X1 port map( A1 => n20509, A2 => n20053, B1 => n3986, B2 => 
                           n20058, ZN => n8546);
   U6064 : OAI22_X1 port map( A1 => n20512, A2 => n20054, B1 => n3985, B2 => 
                           n20057, ZN => n8547);
   U6065 : OAI22_X1 port map( A1 => n20515, A2 => n20053, B1 => n3984, B2 => 
                           n20057, ZN => n8548);
   U6066 : OAI22_X1 port map( A1 => n20518, A2 => n20052, B1 => n3983, B2 => 
                           n20057, ZN => n8549);
   U6067 : OAI22_X1 port map( A1 => n20521, A2 => n20052, B1 => n3982, B2 => 
                           n20057, ZN => n8550);
   U6068 : OAI22_X1 port map( A1 => n20524, A2 => n20054, B1 => n3981, B2 => 
                           n20056, ZN => n8551);
   U6069 : OAI22_X1 port map( A1 => n20527, A2 => n20053, B1 => n3980, B2 => 
                           n20056, ZN => n8552);
   U6070 : OAI22_X1 port map( A1 => n20530, A2 => n20052, B1 => n3979, B2 => 
                           n20056, ZN => n8553);
   U6071 : OAI22_X1 port map( A1 => n20533, A2 => n20054, B1 => n3978, B2 => 
                           n20056, ZN => n8554);
   U6072 : OAI22_X1 port map( A1 => n20536, A2 => n20054, B1 => n3977, B2 => 
                           n20055, ZN => n8555);
   U6073 : OAI22_X1 port map( A1 => n20539, A2 => n20053, B1 => n3976, B2 => 
                           n20055, ZN => n8556);
   U6074 : OAI22_X1 port map( A1 => n20542, A2 => n20052, B1 => n3975, B2 => 
                           n20055, ZN => n8557);
   U6075 : OAI22_X1 port map( A1 => n20573, A2 => n20053, B1 => n3974, B2 => 
                           n20055, ZN => n8558);
   U6076 : OAI22_X1 port map( A1 => n20368, A2 => n19942, B1 => n4305, B2 => 
                           n19957, ZN => n8243);
   U6077 : OAI22_X1 port map( A1 => n20371, A2 => n19942, B1 => n4304, B2 => 
                           n19957, ZN => n8244);
   U6078 : OAI22_X1 port map( A1 => n20374, A2 => n19942, B1 => n4303, B2 => 
                           n19957, ZN => n8245);
   U6079 : OAI22_X1 port map( A1 => n20377, A2 => n19942, B1 => n4302, B2 => 
                           n19957, ZN => n8246);
   U6080 : OAI22_X1 port map( A1 => n20380, A2 => n19942, B1 => n4301, B2 => 
                           n19956, ZN => n8247);
   U6081 : OAI22_X1 port map( A1 => n20383, A2 => n19942, B1 => n4300, B2 => 
                           n19956, ZN => n8248);
   U6082 : OAI22_X1 port map( A1 => n20386, A2 => n19942, B1 => n4299, B2 => 
                           n19956, ZN => n8249);
   U6083 : OAI22_X1 port map( A1 => n20389, A2 => n19942, B1 => n4298, B2 => 
                           n19956, ZN => n8250);
   U6084 : OAI22_X1 port map( A1 => n20392, A2 => n19942, B1 => n4297, B2 => 
                           n19955, ZN => n8251);
   U6085 : OAI22_X1 port map( A1 => n20395, A2 => n19942, B1 => n4296, B2 => 
                           n19955, ZN => n8252);
   U6086 : OAI22_X1 port map( A1 => n20398, A2 => n19942, B1 => n4295, B2 => 
                           n19955, ZN => n8253);
   U6087 : OAI22_X1 port map( A1 => n20401, A2 => n19942, B1 => n4294, B2 => 
                           n19955, ZN => n8254);
   U6088 : OAI22_X1 port map( A1 => n20404, A2 => n19941, B1 => n4293, B2 => 
                           n19954, ZN => n8255);
   U6089 : OAI22_X1 port map( A1 => n20407, A2 => n19941, B1 => n4292, B2 => 
                           n19954, ZN => n8256);
   U6090 : OAI22_X1 port map( A1 => n20410, A2 => n19941, B1 => n4291, B2 => 
                           n19954, ZN => n8257);
   U6091 : OAI22_X1 port map( A1 => n20413, A2 => n19941, B1 => n4290, B2 => 
                           n19954, ZN => n8258);
   U6092 : OAI22_X1 port map( A1 => n20416, A2 => n19941, B1 => n4289, B2 => 
                           n19953, ZN => n8259);
   U6093 : OAI22_X1 port map( A1 => n20419, A2 => n19941, B1 => n4288, B2 => 
                           n19953, ZN => n8260);
   U6094 : OAI22_X1 port map( A1 => n20422, A2 => n19941, B1 => n4287, B2 => 
                           n19953, ZN => n8261);
   U6095 : OAI22_X1 port map( A1 => n20425, A2 => n19941, B1 => n4286, B2 => 
                           n19953, ZN => n8262);
   U6096 : OAI22_X1 port map( A1 => n20428, A2 => n19941, B1 => n4285, B2 => 
                           n19952, ZN => n8263);
   U6097 : OAI22_X1 port map( A1 => n20431, A2 => n19941, B1 => n4284, B2 => 
                           n19952, ZN => n8264);
   U6098 : OAI22_X1 port map( A1 => n20434, A2 => n19941, B1 => n4283, B2 => 
                           n19952, ZN => n8265);
   U6099 : OAI22_X1 port map( A1 => n20437, A2 => n19941, B1 => n4282, B2 => 
                           n19952, ZN => n8266);
   U6100 : OAI22_X1 port map( A1 => n20440, A2 => n19940, B1 => n4281, B2 => 
                           n19951, ZN => n8267);
   U6101 : OAI22_X1 port map( A1 => n20443, A2 => n19940, B1 => n4280, B2 => 
                           n19951, ZN => n8268);
   U6102 : OAI22_X1 port map( A1 => n20446, A2 => n19940, B1 => n4279, B2 => 
                           n19951, ZN => n8269);
   U6103 : OAI22_X1 port map( A1 => n20449, A2 => n19940, B1 => n4278, B2 => 
                           n19951, ZN => n8270);
   U6104 : OAI22_X1 port map( A1 => n20452, A2 => n19940, B1 => n4277, B2 => 
                           n19950, ZN => n8271);
   U6105 : OAI22_X1 port map( A1 => n20455, A2 => n19940, B1 => n4276, B2 => 
                           n19950, ZN => n8272);
   U6106 : OAI22_X1 port map( A1 => n20458, A2 => n19940, B1 => n4275, B2 => 
                           n19950, ZN => n8273);
   U6107 : OAI22_X1 port map( A1 => n20461, A2 => n19940, B1 => n4274, B2 => 
                           n19950, ZN => n8274);
   U6108 : OAI22_X1 port map( A1 => n20464, A2 => n19940, B1 => n4273, B2 => 
                           n19949, ZN => n8275);
   U6109 : OAI22_X1 port map( A1 => n20467, A2 => n19940, B1 => n4272, B2 => 
                           n19949, ZN => n8276);
   U6110 : OAI22_X1 port map( A1 => n20470, A2 => n19940, B1 => n4271, B2 => 
                           n19949, ZN => n8277);
   U6111 : OAI22_X1 port map( A1 => n20473, A2 => n19940, B1 => n4270, B2 => 
                           n19949, ZN => n8278);
   U6112 : OAI22_X1 port map( A1 => n20476, A2 => n19942, B1 => n4269, B2 => 
                           n19948, ZN => n8279);
   U6113 : OAI22_X1 port map( A1 => n20479, A2 => n19941, B1 => n4268, B2 => 
                           n19948, ZN => n8280);
   U6114 : OAI22_X1 port map( A1 => n20482, A2 => n19940, B1 => n4267, B2 => 
                           n19948, ZN => n8281);
   U6115 : OAI22_X1 port map( A1 => n20485, A2 => n19942, B1 => n4266, B2 => 
                           n19948, ZN => n8282);
   U6116 : OAI22_X1 port map( A1 => n20488, A2 => n19941, B1 => n4265, B2 => 
                           n19947, ZN => n8283);
   U6117 : OAI22_X1 port map( A1 => n20491, A2 => n19940, B1 => n4264, B2 => 
                           n19947, ZN => n8284);
   U6118 : OAI22_X1 port map( A1 => n20494, A2 => n19942, B1 => n4263, B2 => 
                           n19947, ZN => n8285);
   U6119 : OAI22_X1 port map( A1 => n20497, A2 => n19941, B1 => n4262, B2 => 
                           n19947, ZN => n8286);
   U6120 : OAI22_X1 port map( A1 => n20500, A2 => n19940, B1 => n4261, B2 => 
                           n19946, ZN => n8287);
   U6121 : OAI22_X1 port map( A1 => n20503, A2 => n19942, B1 => n4260, B2 => 
                           n19946, ZN => n8288);
   U6122 : OAI22_X1 port map( A1 => n20506, A2 => n19941, B1 => n4259, B2 => 
                           n19946, ZN => n8289);
   U6123 : OAI22_X1 port map( A1 => n20509, A2 => n19941, B1 => n4258, B2 => 
                           n19946, ZN => n8290);
   U6124 : OAI22_X1 port map( A1 => n20512, A2 => n19942, B1 => n4257, B2 => 
                           n19945, ZN => n8291);
   U6125 : OAI22_X1 port map( A1 => n20515, A2 => n19941, B1 => n4256, B2 => 
                           n19945, ZN => n8292);
   U6126 : OAI22_X1 port map( A1 => n20518, A2 => n19940, B1 => n4255, B2 => 
                           n19945, ZN => n8293);
   U6127 : OAI22_X1 port map( A1 => n20521, A2 => n19940, B1 => n4254, B2 => 
                           n19945, ZN => n8294);
   U6128 : OAI22_X1 port map( A1 => n20524, A2 => n19942, B1 => n4253, B2 => 
                           n19944, ZN => n8295);
   U6129 : OAI22_X1 port map( A1 => n20527, A2 => n19941, B1 => n4252, B2 => 
                           n19944, ZN => n8296);
   U6130 : OAI22_X1 port map( A1 => n20530, A2 => n19940, B1 => n4251, B2 => 
                           n19944, ZN => n8297);
   U6131 : OAI22_X1 port map( A1 => n20533, A2 => n19942, B1 => n4250, B2 => 
                           n19944, ZN => n8298);
   U6132 : OAI22_X1 port map( A1 => n20536, A2 => n19942, B1 => n4249, B2 => 
                           n19943, ZN => n8299);
   U6133 : OAI22_X1 port map( A1 => n20539, A2 => n19941, B1 => n4248, B2 => 
                           n19943, ZN => n8300);
   U6134 : OAI22_X1 port map( A1 => n20542, A2 => n19940, B1 => n4247, B2 => 
                           n19943, ZN => n8301);
   U6135 : OAI22_X1 port map( A1 => n20573, A2 => n19941, B1 => n4246, B2 => 
                           n19943, ZN => n8302);
   U6136 : OAI22_X1 port map( A1 => n20369, A2 => n20194, B1 => n3700, B2 => 
                           n20209, ZN => n8819);
   U6137 : OAI22_X1 port map( A1 => n20372, A2 => n20194, B1 => n3699, B2 => 
                           n20209, ZN => n8820);
   U6138 : OAI22_X1 port map( A1 => n20375, A2 => n20194, B1 => n3698, B2 => 
                           n20209, ZN => n8821);
   U6139 : OAI22_X1 port map( A1 => n20378, A2 => n20194, B1 => n3697, B2 => 
                           n20209, ZN => n8822);
   U6140 : OAI22_X1 port map( A1 => n20381, A2 => n20194, B1 => n3696, B2 => 
                           n20208, ZN => n8823);
   U6141 : OAI22_X1 port map( A1 => n20384, A2 => n20194, B1 => n3695, B2 => 
                           n20208, ZN => n8824);
   U6142 : OAI22_X1 port map( A1 => n20387, A2 => n20194, B1 => n3694, B2 => 
                           n20208, ZN => n8825);
   U6143 : OAI22_X1 port map( A1 => n20390, A2 => n20194, B1 => n3693, B2 => 
                           n20208, ZN => n8826);
   U6144 : OAI22_X1 port map( A1 => n20393, A2 => n20194, B1 => n3692, B2 => 
                           n20207, ZN => n8827);
   U6145 : OAI22_X1 port map( A1 => n20396, A2 => n20194, B1 => n3691, B2 => 
                           n20207, ZN => n8828);
   U6146 : OAI22_X1 port map( A1 => n20399, A2 => n20194, B1 => n3690, B2 => 
                           n20207, ZN => n8829);
   U6147 : OAI22_X1 port map( A1 => n20402, A2 => n20194, B1 => n3689, B2 => 
                           n20207, ZN => n8830);
   U6148 : OAI22_X1 port map( A1 => n20405, A2 => n20193, B1 => n3688, B2 => 
                           n20206, ZN => n8831);
   U6149 : OAI22_X1 port map( A1 => n20408, A2 => n20193, B1 => n3687, B2 => 
                           n20206, ZN => n8832);
   U6150 : OAI22_X1 port map( A1 => n20411, A2 => n20193, B1 => n3686, B2 => 
                           n20206, ZN => n8833);
   U6151 : OAI22_X1 port map( A1 => n20414, A2 => n20193, B1 => n3685, B2 => 
                           n20206, ZN => n8834);
   U6152 : OAI22_X1 port map( A1 => n20417, A2 => n20193, B1 => n3684, B2 => 
                           n20205, ZN => n8835);
   U6153 : OAI22_X1 port map( A1 => n20420, A2 => n20193, B1 => n3683, B2 => 
                           n20205, ZN => n8836);
   U6154 : OAI22_X1 port map( A1 => n20423, A2 => n20193, B1 => n3682, B2 => 
                           n20205, ZN => n8837);
   U6155 : OAI22_X1 port map( A1 => n20426, A2 => n20193, B1 => n3681, B2 => 
                           n20205, ZN => n8838);
   U6156 : OAI22_X1 port map( A1 => n20429, A2 => n20193, B1 => n3680, B2 => 
                           n20204, ZN => n8839);
   U6157 : OAI22_X1 port map( A1 => n20432, A2 => n20193, B1 => n3679, B2 => 
                           n20204, ZN => n8840);
   U6158 : OAI22_X1 port map( A1 => n20435, A2 => n20193, B1 => n3678, B2 => 
                           n20204, ZN => n8841);
   U6159 : OAI22_X1 port map( A1 => n20438, A2 => n20193, B1 => n3677, B2 => 
                           n20204, ZN => n8842);
   U6160 : OAI22_X1 port map( A1 => n20441, A2 => n20192, B1 => n3676, B2 => 
                           n20203, ZN => n8843);
   U6161 : OAI22_X1 port map( A1 => n20444, A2 => n20192, B1 => n3675, B2 => 
                           n20203, ZN => n8844);
   U6162 : OAI22_X1 port map( A1 => n20447, A2 => n20192, B1 => n3674, B2 => 
                           n20203, ZN => n8845);
   U6163 : OAI22_X1 port map( A1 => n20450, A2 => n20192, B1 => n3673, B2 => 
                           n20203, ZN => n8846);
   U6164 : OAI22_X1 port map( A1 => n20453, A2 => n20192, B1 => n3672, B2 => 
                           n20202, ZN => n8847);
   U6165 : OAI22_X1 port map( A1 => n20456, A2 => n20192, B1 => n3671, B2 => 
                           n20202, ZN => n8848);
   U6166 : OAI22_X1 port map( A1 => n20459, A2 => n20192, B1 => n3670, B2 => 
                           n20202, ZN => n8849);
   U6167 : OAI22_X1 port map( A1 => n20462, A2 => n20192, B1 => n3669, B2 => 
                           n20202, ZN => n8850);
   U6168 : OAI22_X1 port map( A1 => n20465, A2 => n20192, B1 => n3668, B2 => 
                           n20201, ZN => n8851);
   U6169 : OAI22_X1 port map( A1 => n20468, A2 => n20192, B1 => n3667, B2 => 
                           n20201, ZN => n8852);
   U6170 : OAI22_X1 port map( A1 => n20471, A2 => n20192, B1 => n3666, B2 => 
                           n20201, ZN => n8853);
   U6171 : OAI22_X1 port map( A1 => n20474, A2 => n20192, B1 => n3665, B2 => 
                           n20201, ZN => n8854);
   U6172 : OAI22_X1 port map( A1 => n20477, A2 => n20194, B1 => n3664, B2 => 
                           n20200, ZN => n8855);
   U6173 : OAI22_X1 port map( A1 => n20480, A2 => n20193, B1 => n3663, B2 => 
                           n20200, ZN => n8856);
   U6174 : OAI22_X1 port map( A1 => n20483, A2 => n20192, B1 => n3662, B2 => 
                           n20200, ZN => n8857);
   U6175 : OAI22_X1 port map( A1 => n20486, A2 => n20194, B1 => n3661, B2 => 
                           n20200, ZN => n8858);
   U6176 : OAI22_X1 port map( A1 => n20489, A2 => n20193, B1 => n3660, B2 => 
                           n20199, ZN => n8859);
   U6177 : OAI22_X1 port map( A1 => n20492, A2 => n20192, B1 => n3659, B2 => 
                           n20199, ZN => n8860);
   U6178 : OAI22_X1 port map( A1 => n20495, A2 => n20194, B1 => n3658, B2 => 
                           n20199, ZN => n8861);
   U6179 : OAI22_X1 port map( A1 => n20498, A2 => n20193, B1 => n3657, B2 => 
                           n20199, ZN => n8862);
   U6180 : OAI22_X1 port map( A1 => n20501, A2 => n20192, B1 => n3656, B2 => 
                           n20198, ZN => n8863);
   U6181 : OAI22_X1 port map( A1 => n20504, A2 => n20194, B1 => n3655, B2 => 
                           n20198, ZN => n8864);
   U6182 : OAI22_X1 port map( A1 => n20507, A2 => n20193, B1 => n3654, B2 => 
                           n20198, ZN => n8865);
   U6183 : OAI22_X1 port map( A1 => n20510, A2 => n20193, B1 => n3653, B2 => 
                           n20198, ZN => n8866);
   U6184 : OAI22_X1 port map( A1 => n20513, A2 => n20194, B1 => n3652, B2 => 
                           n20197, ZN => n8867);
   U6185 : OAI22_X1 port map( A1 => n20516, A2 => n20193, B1 => n3651, B2 => 
                           n20197, ZN => n8868);
   U6186 : OAI22_X1 port map( A1 => n20519, A2 => n20192, B1 => n3650, B2 => 
                           n20197, ZN => n8869);
   U6187 : OAI22_X1 port map( A1 => n20522, A2 => n20192, B1 => n3649, B2 => 
                           n20197, ZN => n8870);
   U6188 : OAI22_X1 port map( A1 => n20525, A2 => n20194, B1 => n3648, B2 => 
                           n20196, ZN => n8871);
   U6189 : OAI22_X1 port map( A1 => n20528, A2 => n20193, B1 => n3647, B2 => 
                           n20196, ZN => n8872);
   U6190 : OAI22_X1 port map( A1 => n20531, A2 => n20192, B1 => n3646, B2 => 
                           n20196, ZN => n8873);
   U6191 : OAI22_X1 port map( A1 => n20534, A2 => n20194, B1 => n3645, B2 => 
                           n20196, ZN => n8874);
   U6192 : OAI22_X1 port map( A1 => n20537, A2 => n20194, B1 => n3644, B2 => 
                           n20195, ZN => n8875);
   U6193 : OAI22_X1 port map( A1 => n20540, A2 => n20193, B1 => n3643, B2 => 
                           n20195, ZN => n8876);
   U6194 : OAI22_X1 port map( A1 => n20543, A2 => n20192, B1 => n3642, B2 => 
                           n20195, ZN => n8877);
   U6195 : OAI22_X1 port map( A1 => n20574, A2 => n20193, B1 => n3641, B2 => 
                           n20195, ZN => n8878);
   U6196 : OAI22_X1 port map( A1 => n20356, A2 => n20053, B1 => n4037, B2 => 
                           n20070, ZN => n8495);
   U6197 : OAI22_X1 port map( A1 => n20359, A2 => n20052, B1 => n4036, B2 => 
                           n20070, ZN => n8496);
   U6198 : OAI22_X1 port map( A1 => n20362, A2 => n20052, B1 => n4035, B2 => 
                           n20070, ZN => n8497);
   U6199 : OAI22_X1 port map( A1 => n20365, A2 => n20054, B1 => n4034, B2 => 
                           n20070, ZN => n8498);
   U6200 : OAI22_X1 port map( A1 => n20356, A2 => n19941, B1 => n4309, B2 => 
                           n19958, ZN => n8239);
   U6201 : OAI22_X1 port map( A1 => n20359, A2 => n19940, B1 => n4308, B2 => 
                           n19958, ZN => n8240);
   U6202 : OAI22_X1 port map( A1 => n20362, A2 => n19940, B1 => n4307, B2 => 
                           n19958, ZN => n8241);
   U6203 : OAI22_X1 port map( A1 => n20365, A2 => n19942, B1 => n4306, B2 => 
                           n19958, ZN => n8242);
   U6204 : OAI22_X1 port map( A1 => n20357, A2 => n20193, B1 => n3704, B2 => 
                           n20210, ZN => n8815);
   U6205 : OAI22_X1 port map( A1 => n20360, A2 => n20192, B1 => n3703, B2 => 
                           n20210, ZN => n8816);
   U6206 : OAI22_X1 port map( A1 => n20363, A2 => n20192, B1 => n3702, B2 => 
                           n20210, ZN => n8817);
   U6207 : OAI22_X1 port map( A1 => n20366, A2 => n20194, B1 => n3701, B2 => 
                           n20210, ZN => n8818);
   U6208 : OAI22_X1 port map( A1 => n20368, A2 => n20026, B1 => n4099, B2 => 
                           n20041, ZN => n8435);
   U6209 : OAI22_X1 port map( A1 => n20371, A2 => n20026, B1 => n4098, B2 => 
                           n20041, ZN => n8436);
   U6210 : OAI22_X1 port map( A1 => n20374, A2 => n20026, B1 => n4097, B2 => 
                           n20041, ZN => n8437);
   U6211 : OAI22_X1 port map( A1 => n20377, A2 => n20026, B1 => n4096, B2 => 
                           n20041, ZN => n8438);
   U6212 : OAI22_X1 port map( A1 => n20380, A2 => n20026, B1 => n4095, B2 => 
                           n20040, ZN => n8439);
   U6213 : OAI22_X1 port map( A1 => n20383, A2 => n20026, B1 => n4094, B2 => 
                           n20040, ZN => n8440);
   U6214 : OAI22_X1 port map( A1 => n20386, A2 => n20026, B1 => n4093, B2 => 
                           n20040, ZN => n8441);
   U6215 : OAI22_X1 port map( A1 => n20389, A2 => n20026, B1 => n4092, B2 => 
                           n20040, ZN => n8442);
   U6216 : OAI22_X1 port map( A1 => n20392, A2 => n20026, B1 => n4091, B2 => 
                           n20039, ZN => n8443);
   U6217 : OAI22_X1 port map( A1 => n20395, A2 => n20026, B1 => n4090, B2 => 
                           n20039, ZN => n8444);
   U6218 : OAI22_X1 port map( A1 => n20398, A2 => n20026, B1 => n4089, B2 => 
                           n20039, ZN => n8445);
   U6219 : OAI22_X1 port map( A1 => n20401, A2 => n20026, B1 => n4088, B2 => 
                           n20039, ZN => n8446);
   U6220 : OAI22_X1 port map( A1 => n20404, A2 => n20025, B1 => n4087, B2 => 
                           n20038, ZN => n8447);
   U6221 : OAI22_X1 port map( A1 => n20407, A2 => n20025, B1 => n4086, B2 => 
                           n20038, ZN => n8448);
   U6222 : OAI22_X1 port map( A1 => n20410, A2 => n20025, B1 => n4085, B2 => 
                           n20038, ZN => n8449);
   U6223 : OAI22_X1 port map( A1 => n20413, A2 => n20025, B1 => n4084, B2 => 
                           n20038, ZN => n8450);
   U6224 : OAI22_X1 port map( A1 => n20416, A2 => n20025, B1 => n4083, B2 => 
                           n20037, ZN => n8451);
   U6225 : OAI22_X1 port map( A1 => n20419, A2 => n20025, B1 => n4082, B2 => 
                           n20037, ZN => n8452);
   U6226 : OAI22_X1 port map( A1 => n20422, A2 => n20025, B1 => n4081, B2 => 
                           n20037, ZN => n8453);
   U6227 : OAI22_X1 port map( A1 => n20425, A2 => n20025, B1 => n4080, B2 => 
                           n20037, ZN => n8454);
   U6228 : OAI22_X1 port map( A1 => n20428, A2 => n20025, B1 => n4079, B2 => 
                           n20036, ZN => n8455);
   U6229 : OAI22_X1 port map( A1 => n20431, A2 => n20025, B1 => n4078, B2 => 
                           n20036, ZN => n8456);
   U6230 : OAI22_X1 port map( A1 => n20434, A2 => n20025, B1 => n4077, B2 => 
                           n20036, ZN => n8457);
   U6231 : OAI22_X1 port map( A1 => n20437, A2 => n20025, B1 => n4076, B2 => 
                           n20036, ZN => n8458);
   U6232 : OAI22_X1 port map( A1 => n20440, A2 => n20024, B1 => n4075, B2 => 
                           n20035, ZN => n8459);
   U6233 : OAI22_X1 port map( A1 => n20443, A2 => n20024, B1 => n4074, B2 => 
                           n20035, ZN => n8460);
   U6234 : OAI22_X1 port map( A1 => n20446, A2 => n20024, B1 => n4073, B2 => 
                           n20035, ZN => n8461);
   U6235 : OAI22_X1 port map( A1 => n20449, A2 => n20024, B1 => n4072, B2 => 
                           n20035, ZN => n8462);
   U6236 : OAI22_X1 port map( A1 => n20452, A2 => n20024, B1 => n4071, B2 => 
                           n20034, ZN => n8463);
   U6237 : OAI22_X1 port map( A1 => n20455, A2 => n20024, B1 => n4070, B2 => 
                           n20034, ZN => n8464);
   U6238 : OAI22_X1 port map( A1 => n20458, A2 => n20024, B1 => n4069, B2 => 
                           n20034, ZN => n8465);
   U6239 : OAI22_X1 port map( A1 => n20461, A2 => n20024, B1 => n4068, B2 => 
                           n20034, ZN => n8466);
   U6240 : OAI22_X1 port map( A1 => n20464, A2 => n20024, B1 => n4067, B2 => 
                           n20033, ZN => n8467);
   U6241 : OAI22_X1 port map( A1 => n20467, A2 => n20024, B1 => n4066, B2 => 
                           n20033, ZN => n8468);
   U6242 : OAI22_X1 port map( A1 => n20470, A2 => n20024, B1 => n4065, B2 => 
                           n20033, ZN => n8469);
   U6243 : OAI22_X1 port map( A1 => n20473, A2 => n20024, B1 => n4064, B2 => 
                           n20033, ZN => n8470);
   U6244 : OAI22_X1 port map( A1 => n20476, A2 => n20026, B1 => n4063, B2 => 
                           n20032, ZN => n8471);
   U6245 : OAI22_X1 port map( A1 => n20479, A2 => n20025, B1 => n4062, B2 => 
                           n20032, ZN => n8472);
   U6246 : OAI22_X1 port map( A1 => n20482, A2 => n20024, B1 => n4061, B2 => 
                           n20032, ZN => n8473);
   U6247 : OAI22_X1 port map( A1 => n20485, A2 => n20026, B1 => n4060, B2 => 
                           n20032, ZN => n8474);
   U6248 : OAI22_X1 port map( A1 => n20488, A2 => n20025, B1 => n4059, B2 => 
                           n20031, ZN => n8475);
   U6249 : OAI22_X1 port map( A1 => n20491, A2 => n20024, B1 => n4058, B2 => 
                           n20031, ZN => n8476);
   U6250 : OAI22_X1 port map( A1 => n20494, A2 => n20026, B1 => n4057, B2 => 
                           n20031, ZN => n8477);
   U6251 : OAI22_X1 port map( A1 => n20497, A2 => n20025, B1 => n4056, B2 => 
                           n20031, ZN => n8478);
   U6252 : OAI22_X1 port map( A1 => n20500, A2 => n20024, B1 => n4055, B2 => 
                           n20030, ZN => n8479);
   U6253 : OAI22_X1 port map( A1 => n20503, A2 => n20026, B1 => n4054, B2 => 
                           n20030, ZN => n8480);
   U6254 : OAI22_X1 port map( A1 => n20506, A2 => n20025, B1 => n4053, B2 => 
                           n20030, ZN => n8481);
   U6255 : OAI22_X1 port map( A1 => n20509, A2 => n20025, B1 => n4052, B2 => 
                           n20030, ZN => n8482);
   U6256 : OAI22_X1 port map( A1 => n20512, A2 => n20026, B1 => n4051, B2 => 
                           n20029, ZN => n8483);
   U6257 : OAI22_X1 port map( A1 => n20515, A2 => n20025, B1 => n4050, B2 => 
                           n20029, ZN => n8484);
   U6258 : OAI22_X1 port map( A1 => n20518, A2 => n20024, B1 => n4049, B2 => 
                           n20029, ZN => n8485);
   U6259 : OAI22_X1 port map( A1 => n20521, A2 => n20024, B1 => n4048, B2 => 
                           n20029, ZN => n8486);
   U6260 : OAI22_X1 port map( A1 => n20524, A2 => n20026, B1 => n4047, B2 => 
                           n20028, ZN => n8487);
   U6261 : OAI22_X1 port map( A1 => n20527, A2 => n20025, B1 => n4046, B2 => 
                           n20028, ZN => n8488);
   U6262 : OAI22_X1 port map( A1 => n20530, A2 => n20024, B1 => n4045, B2 => 
                           n20028, ZN => n8489);
   U6263 : OAI22_X1 port map( A1 => n20533, A2 => n20026, B1 => n4044, B2 => 
                           n20028, ZN => n8490);
   U6264 : OAI22_X1 port map( A1 => n20536, A2 => n20026, B1 => n4043, B2 => 
                           n20027, ZN => n8491);
   U6265 : OAI22_X1 port map( A1 => n20539, A2 => n20025, B1 => n4042, B2 => 
                           n20027, ZN => n8492);
   U6266 : OAI22_X1 port map( A1 => n20542, A2 => n20024, B1 => n4041, B2 => 
                           n20027, ZN => n8493);
   U6267 : OAI22_X1 port map( A1 => n20573, A2 => n20025, B1 => n4040, B2 => 
                           n20027, ZN => n8494);
   U6268 : OAI22_X1 port map( A1 => n20369, A2 => n20554, B1 => n3287, B2 => 
                           n20569, ZN => n9203);
   U6269 : OAI22_X1 port map( A1 => n20372, A2 => n20554, B1 => n3285, B2 => 
                           n20569, ZN => n9204);
   U6270 : OAI22_X1 port map( A1 => n20375, A2 => n20554, B1 => n3283, B2 => 
                           n20569, ZN => n9205);
   U6271 : OAI22_X1 port map( A1 => n20378, A2 => n20554, B1 => n3281, B2 => 
                           n20569, ZN => n9206);
   U6272 : OAI22_X1 port map( A1 => n20381, A2 => n20554, B1 => n3279, B2 => 
                           n20568, ZN => n9207);
   U6273 : OAI22_X1 port map( A1 => n20384, A2 => n20554, B1 => n3277, B2 => 
                           n20568, ZN => n9208);
   U6274 : OAI22_X1 port map( A1 => n20387, A2 => n20554, B1 => n3275, B2 => 
                           n20568, ZN => n9209);
   U6275 : OAI22_X1 port map( A1 => n20390, A2 => n20554, B1 => n3273, B2 => 
                           n20568, ZN => n9210);
   U6276 : OAI22_X1 port map( A1 => n20393, A2 => n20554, B1 => n3271, B2 => 
                           n20567, ZN => n9211);
   U6277 : OAI22_X1 port map( A1 => n20396, A2 => n20554, B1 => n3269, B2 => 
                           n20567, ZN => n9212);
   U6278 : OAI22_X1 port map( A1 => n20399, A2 => n20554, B1 => n3267, B2 => 
                           n20567, ZN => n9213);
   U6279 : OAI22_X1 port map( A1 => n20402, A2 => n20554, B1 => n3265, B2 => 
                           n20567, ZN => n9214);
   U6280 : OAI22_X1 port map( A1 => n20405, A2 => n20553, B1 => n3263, B2 => 
                           n20566, ZN => n9215);
   U6281 : OAI22_X1 port map( A1 => n20408, A2 => n20553, B1 => n3261, B2 => 
                           n20566, ZN => n9216);
   U6282 : OAI22_X1 port map( A1 => n20411, A2 => n20553, B1 => n3259, B2 => 
                           n20566, ZN => n9217);
   U6283 : OAI22_X1 port map( A1 => n20414, A2 => n20553, B1 => n3257, B2 => 
                           n20566, ZN => n9218);
   U6284 : OAI22_X1 port map( A1 => n20417, A2 => n20553, B1 => n3255, B2 => 
                           n20565, ZN => n9219);
   U6285 : OAI22_X1 port map( A1 => n20420, A2 => n20553, B1 => n3253, B2 => 
                           n20565, ZN => n9220);
   U6286 : OAI22_X1 port map( A1 => n20423, A2 => n20553, B1 => n3251, B2 => 
                           n20565, ZN => n9221);
   U6287 : OAI22_X1 port map( A1 => n20426, A2 => n20553, B1 => n3249, B2 => 
                           n20565, ZN => n9222);
   U6288 : OAI22_X1 port map( A1 => n20429, A2 => n20553, B1 => n3247, B2 => 
                           n20564, ZN => n9223);
   U6289 : OAI22_X1 port map( A1 => n20432, A2 => n20553, B1 => n3245, B2 => 
                           n20564, ZN => n9224);
   U6290 : OAI22_X1 port map( A1 => n20435, A2 => n20553, B1 => n3243, B2 => 
                           n20564, ZN => n9225);
   U6291 : OAI22_X1 port map( A1 => n20438, A2 => n20553, B1 => n3241, B2 => 
                           n20564, ZN => n9226);
   U6292 : OAI22_X1 port map( A1 => n20441, A2 => n20552, B1 => n3239, B2 => 
                           n20563, ZN => n9227);
   U6293 : OAI22_X1 port map( A1 => n20444, A2 => n20552, B1 => n3237, B2 => 
                           n20563, ZN => n9228);
   U6294 : OAI22_X1 port map( A1 => n20447, A2 => n20552, B1 => n3235, B2 => 
                           n20563, ZN => n9229);
   U6295 : OAI22_X1 port map( A1 => n20450, A2 => n20552, B1 => n3233, B2 => 
                           n20563, ZN => n9230);
   U6296 : OAI22_X1 port map( A1 => n20453, A2 => n20552, B1 => n3231, B2 => 
                           n20562, ZN => n9231);
   U6297 : OAI22_X1 port map( A1 => n20456, A2 => n20552, B1 => n3229, B2 => 
                           n20562, ZN => n9232);
   U6298 : OAI22_X1 port map( A1 => n20459, A2 => n20552, B1 => n3227, B2 => 
                           n20562, ZN => n9233);
   U6299 : OAI22_X1 port map( A1 => n20462, A2 => n20552, B1 => n3225, B2 => 
                           n20562, ZN => n9234);
   U6300 : OAI22_X1 port map( A1 => n20465, A2 => n20552, B1 => n3223, B2 => 
                           n20561, ZN => n9235);
   U6301 : OAI22_X1 port map( A1 => n20468, A2 => n20552, B1 => n3221, B2 => 
                           n20561, ZN => n9236);
   U6302 : OAI22_X1 port map( A1 => n20471, A2 => n20552, B1 => n3219, B2 => 
                           n20561, ZN => n9237);
   U6303 : OAI22_X1 port map( A1 => n20474, A2 => n20552, B1 => n3217, B2 => 
                           n20561, ZN => n9238);
   U6304 : OAI22_X1 port map( A1 => n20477, A2 => n20554, B1 => n3215, B2 => 
                           n20560, ZN => n9239);
   U6305 : OAI22_X1 port map( A1 => n20480, A2 => n20553, B1 => n3213, B2 => 
                           n20560, ZN => n9240);
   U6306 : OAI22_X1 port map( A1 => n20483, A2 => n20552, B1 => n3211, B2 => 
                           n20560, ZN => n9241);
   U6307 : OAI22_X1 port map( A1 => n20486, A2 => n20554, B1 => n3209, B2 => 
                           n20560, ZN => n9242);
   U6308 : OAI22_X1 port map( A1 => n20489, A2 => n20553, B1 => n3207, B2 => 
                           n20559, ZN => n9243);
   U6309 : OAI22_X1 port map( A1 => n20492, A2 => n20552, B1 => n3205, B2 => 
                           n20559, ZN => n9244);
   U6310 : OAI22_X1 port map( A1 => n20495, A2 => n20554, B1 => n3203, B2 => 
                           n20559, ZN => n9245);
   U6311 : OAI22_X1 port map( A1 => n20498, A2 => n20553, B1 => n3201, B2 => 
                           n20559, ZN => n9246);
   U6312 : OAI22_X1 port map( A1 => n20501, A2 => n20552, B1 => n3199, B2 => 
                           n20558, ZN => n9247);
   U6313 : OAI22_X1 port map( A1 => n20504, A2 => n20554, B1 => n3197, B2 => 
                           n20558, ZN => n9248);
   U6314 : OAI22_X1 port map( A1 => n20507, A2 => n20553, B1 => n3195, B2 => 
                           n20558, ZN => n9249);
   U6315 : OAI22_X1 port map( A1 => n20510, A2 => n20553, B1 => n3193, B2 => 
                           n20558, ZN => n9250);
   U6316 : OAI22_X1 port map( A1 => n20513, A2 => n20554, B1 => n3191, B2 => 
                           n20557, ZN => n9251);
   U6317 : OAI22_X1 port map( A1 => n20516, A2 => n20553, B1 => n3189, B2 => 
                           n20557, ZN => n9252);
   U6318 : OAI22_X1 port map( A1 => n20519, A2 => n20552, B1 => n3187, B2 => 
                           n20557, ZN => n9253);
   U6319 : OAI22_X1 port map( A1 => n20522, A2 => n20552, B1 => n3185, B2 => 
                           n20557, ZN => n9254);
   U6320 : OAI22_X1 port map( A1 => n20525, A2 => n20554, B1 => n3183, B2 => 
                           n20556, ZN => n9255);
   U6321 : OAI22_X1 port map( A1 => n20528, A2 => n20553, B1 => n3181, B2 => 
                           n20556, ZN => n9256);
   U6322 : OAI22_X1 port map( A1 => n20531, A2 => n20552, B1 => n3179, B2 => 
                           n20556, ZN => n9257);
   U6323 : OAI22_X1 port map( A1 => n20534, A2 => n20554, B1 => n3177, B2 => 
                           n20556, ZN => n9258);
   U6324 : OAI22_X1 port map( A1 => n20537, A2 => n20554, B1 => n3175, B2 => 
                           n20555, ZN => n9259);
   U6325 : OAI22_X1 port map( A1 => n20540, A2 => n20553, B1 => n3173, B2 => 
                           n20555, ZN => n9260);
   U6326 : OAI22_X1 port map( A1 => n20543, A2 => n20552, B1 => n3171, B2 => 
                           n20555, ZN => n9261);
   U6327 : OAI22_X1 port map( A1 => n20574, A2 => n20553, B1 => n3169, B2 => 
                           n20555, ZN => n9262);
   U6328 : OAI22_X1 port map( A1 => n20356, A2 => n20025, B1 => n4103, B2 => 
                           n20042, ZN => n8431);
   U6329 : OAI22_X1 port map( A1 => n20359, A2 => n20024, B1 => n4102, B2 => 
                           n20042, ZN => n8432);
   U6330 : OAI22_X1 port map( A1 => n20362, A2 => n20024, B1 => n4101, B2 => 
                           n20042, ZN => n8433);
   U6331 : OAI22_X1 port map( A1 => n20365, A2 => n20026, B1 => n4100, B2 => 
                           n20042, ZN => n8434);
   U6332 : OAI22_X1 port map( A1 => n20357, A2 => n20553, B1 => n3295, B2 => 
                           n20570, ZN => n9199);
   U6333 : OAI22_X1 port map( A1 => n20360, A2 => n20552, B1 => n3293, B2 => 
                           n20570, ZN => n9200);
   U6334 : OAI22_X1 port map( A1 => n20363, A2 => n20552, B1 => n3291, B2 => 
                           n20570, ZN => n9201);
   U6335 : OAI22_X1 port map( A1 => n20366, A2 => n20554, B1 => n3289, B2 => 
                           n20570, ZN => n9202);
   U6336 : OAI22_X1 port map( A1 => n20368, A2 => n19914, B1 => n19929, B2 => 
                           n2009, ZN => n8179);
   U6337 : OAI22_X1 port map( A1 => n20371, A2 => n19914, B1 => n19929, B2 => 
                           n2008, ZN => n8180);
   U6338 : OAI22_X1 port map( A1 => n20374, A2 => n19914, B1 => n19929, B2 => 
                           n2007, ZN => n8181);
   U6339 : OAI22_X1 port map( A1 => n20377, A2 => n19914, B1 => n19929, B2 => 
                           n2006, ZN => n8182);
   U6340 : OAI22_X1 port map( A1 => n20380, A2 => n19914, B1 => n19928, B2 => 
                           n2005, ZN => n8183);
   U6341 : OAI22_X1 port map( A1 => n20383, A2 => n19914, B1 => n19928, B2 => 
                           n2004, ZN => n8184);
   U6342 : OAI22_X1 port map( A1 => n20386, A2 => n19914, B1 => n19928, B2 => 
                           n2003, ZN => n8185);
   U6343 : OAI22_X1 port map( A1 => n20389, A2 => n19914, B1 => n19928, B2 => 
                           n2002, ZN => n8186);
   U6344 : OAI22_X1 port map( A1 => n20392, A2 => n19914, B1 => n19927, B2 => 
                           n2001, ZN => n8187);
   U6345 : OAI22_X1 port map( A1 => n20395, A2 => n19914, B1 => n19927, B2 => 
                           n2000, ZN => n8188);
   U6346 : OAI22_X1 port map( A1 => n20398, A2 => n19914, B1 => n19927, B2 => 
                           n1999, ZN => n8189);
   U6347 : OAI22_X1 port map( A1 => n20401, A2 => n19914, B1 => n19927, B2 => 
                           n1998, ZN => n8190);
   U6348 : OAI22_X1 port map( A1 => n20404, A2 => n19913, B1 => n19926, B2 => 
                           n1997, ZN => n8191);
   U6349 : OAI22_X1 port map( A1 => n20407, A2 => n19913, B1 => n19926, B2 => 
                           n1996, ZN => n8192);
   U6350 : OAI22_X1 port map( A1 => n20410, A2 => n19913, B1 => n19926, B2 => 
                           n1995, ZN => n8193);
   U6351 : OAI22_X1 port map( A1 => n20413, A2 => n19913, B1 => n19926, B2 => 
                           n1994, ZN => n8194);
   U6352 : OAI22_X1 port map( A1 => n20416, A2 => n19913, B1 => n19925, B2 => 
                           n1993, ZN => n8195);
   U6353 : OAI22_X1 port map( A1 => n20419, A2 => n19913, B1 => n19925, B2 => 
                           n1992, ZN => n8196);
   U6354 : OAI22_X1 port map( A1 => n20422, A2 => n19913, B1 => n19925, B2 => 
                           n1991, ZN => n8197);
   U6355 : OAI22_X1 port map( A1 => n20425, A2 => n19913, B1 => n19925, B2 => 
                           n1990, ZN => n8198);
   U6356 : OAI22_X1 port map( A1 => n20428, A2 => n19913, B1 => n19924, B2 => 
                           n1989, ZN => n8199);
   U6357 : OAI22_X1 port map( A1 => n20431, A2 => n19913, B1 => n19924, B2 => 
                           n1988, ZN => n8200);
   U6358 : OAI22_X1 port map( A1 => n20434, A2 => n19913, B1 => n19924, B2 => 
                           n1987, ZN => n8201);
   U6359 : OAI22_X1 port map( A1 => n20437, A2 => n19913, B1 => n19924, B2 => 
                           n1986, ZN => n8202);
   U6360 : OAI22_X1 port map( A1 => n20440, A2 => n19912, B1 => n19923, B2 => 
                           n1985, ZN => n8203);
   U6361 : OAI22_X1 port map( A1 => n20443, A2 => n19912, B1 => n19923, B2 => 
                           n1984, ZN => n8204);
   U6362 : OAI22_X1 port map( A1 => n20446, A2 => n19912, B1 => n19923, B2 => 
                           n1983, ZN => n8205);
   U6363 : OAI22_X1 port map( A1 => n20449, A2 => n19912, B1 => n19923, B2 => 
                           n1982, ZN => n8206);
   U6364 : OAI22_X1 port map( A1 => n20452, A2 => n19912, B1 => n19922, B2 => 
                           n1981, ZN => n8207);
   U6365 : OAI22_X1 port map( A1 => n20455, A2 => n19912, B1 => n19922, B2 => 
                           n1980, ZN => n8208);
   U6366 : OAI22_X1 port map( A1 => n20458, A2 => n19912, B1 => n19922, B2 => 
                           n1979, ZN => n8209);
   U6367 : OAI22_X1 port map( A1 => n20461, A2 => n19912, B1 => n19922, B2 => 
                           n1978, ZN => n8210);
   U6368 : OAI22_X1 port map( A1 => n20464, A2 => n19912, B1 => n19921, B2 => 
                           n1977, ZN => n8211);
   U6369 : OAI22_X1 port map( A1 => n20467, A2 => n19912, B1 => n19921, B2 => 
                           n1976, ZN => n8212);
   U6370 : OAI22_X1 port map( A1 => n20470, A2 => n19912, B1 => n19921, B2 => 
                           n1975, ZN => n8213);
   U6371 : OAI22_X1 port map( A1 => n20473, A2 => n19912, B1 => n19921, B2 => 
                           n1974, ZN => n8214);
   U6372 : OAI22_X1 port map( A1 => n20476, A2 => n19914, B1 => n19920, B2 => 
                           n1973, ZN => n8215);
   U6373 : OAI22_X1 port map( A1 => n20479, A2 => n19913, B1 => n19920, B2 => 
                           n1972, ZN => n8216);
   U6374 : OAI22_X1 port map( A1 => n20482, A2 => n19912, B1 => n19920, B2 => 
                           n1971, ZN => n8217);
   U6375 : OAI22_X1 port map( A1 => n20485, A2 => n19914, B1 => n19920, B2 => 
                           n1970, ZN => n8218);
   U6376 : OAI22_X1 port map( A1 => n20488, A2 => n19913, B1 => n19919, B2 => 
                           n1969, ZN => n8219);
   U6377 : OAI22_X1 port map( A1 => n20491, A2 => n19912, B1 => n19919, B2 => 
                           n1968, ZN => n8220);
   U6378 : OAI22_X1 port map( A1 => n20494, A2 => n19914, B1 => n19919, B2 => 
                           n1967, ZN => n8221);
   U6379 : OAI22_X1 port map( A1 => n20497, A2 => n19913, B1 => n19919, B2 => 
                           n1966, ZN => n8222);
   U6380 : OAI22_X1 port map( A1 => n20500, A2 => n19912, B1 => n19918, B2 => 
                           n1965, ZN => n8223);
   U6381 : OAI22_X1 port map( A1 => n20503, A2 => n19914, B1 => n19918, B2 => 
                           n1964, ZN => n8224);
   U6382 : OAI22_X1 port map( A1 => n20506, A2 => n19913, B1 => n19918, B2 => 
                           n1963, ZN => n8225);
   U6383 : OAI22_X1 port map( A1 => n20509, A2 => n19913, B1 => n19918, B2 => 
                           n1962, ZN => n8226);
   U6384 : OAI22_X1 port map( A1 => n20512, A2 => n19914, B1 => n19917, B2 => 
                           n1961, ZN => n8227);
   U6385 : OAI22_X1 port map( A1 => n20515, A2 => n19913, B1 => n19917, B2 => 
                           n1960, ZN => n8228);
   U6386 : OAI22_X1 port map( A1 => n20518, A2 => n19912, B1 => n19917, B2 => 
                           n1959, ZN => n8229);
   U6387 : OAI22_X1 port map( A1 => n20521, A2 => n19912, B1 => n19917, B2 => 
                           n1958, ZN => n8230);
   U6388 : OAI22_X1 port map( A1 => n20524, A2 => n19914, B1 => n19916, B2 => 
                           n1957, ZN => n8231);
   U6389 : OAI22_X1 port map( A1 => n20527, A2 => n19913, B1 => n19916, B2 => 
                           n1956, ZN => n8232);
   U6390 : OAI22_X1 port map( A1 => n20530, A2 => n19912, B1 => n19916, B2 => 
                           n1955, ZN => n8233);
   U6391 : OAI22_X1 port map( A1 => n20533, A2 => n19914, B1 => n19916, B2 => 
                           n1954, ZN => n8234);
   U6392 : OAI22_X1 port map( A1 => n20536, A2 => n19914, B1 => n19915, B2 => 
                           n1953, ZN => n8235);
   U6393 : OAI22_X1 port map( A1 => n20539, A2 => n19913, B1 => n19915, B2 => 
                           n1952, ZN => n8236);
   U6394 : OAI22_X1 port map( A1 => n20542, A2 => n19912, B1 => n19915, B2 => 
                           n1951, ZN => n8237);
   U6395 : OAI22_X1 port map( A1 => n20573, A2 => n19913, B1 => n19915, B2 => 
                           n1950, ZN => n8238);
   U6396 : OAI22_X1 port map( A1 => n20367, A2 => n19606, B1 => n19621, B2 => 
                           n2370, ZN => n7475);
   U6397 : OAI22_X1 port map( A1 => n20370, A2 => n19606, B1 => n19621, B2 => 
                           n2369, ZN => n7476);
   U6398 : OAI22_X1 port map( A1 => n20373, A2 => n19606, B1 => n19621, B2 => 
                           n2368, ZN => n7477);
   U6399 : OAI22_X1 port map( A1 => n20376, A2 => n19606, B1 => n19621, B2 => 
                           n2367, ZN => n7478);
   U6400 : OAI22_X1 port map( A1 => n20379, A2 => n19606, B1 => n19620, B2 => 
                           n2366, ZN => n7479);
   U6401 : OAI22_X1 port map( A1 => n20382, A2 => n19606, B1 => n19620, B2 => 
                           n2365, ZN => n7480);
   U6402 : OAI22_X1 port map( A1 => n20385, A2 => n19606, B1 => n19620, B2 => 
                           n2364, ZN => n7481);
   U6403 : OAI22_X1 port map( A1 => n20388, A2 => n19606, B1 => n19620, B2 => 
                           n2363, ZN => n7482);
   U6404 : OAI22_X1 port map( A1 => n20391, A2 => n19606, B1 => n19619, B2 => 
                           n2362, ZN => n7483);
   U6405 : OAI22_X1 port map( A1 => n20394, A2 => n19606, B1 => n19619, B2 => 
                           n2361, ZN => n7484);
   U6406 : OAI22_X1 port map( A1 => n20397, A2 => n19606, B1 => n19619, B2 => 
                           n2360, ZN => n7485);
   U6407 : OAI22_X1 port map( A1 => n20400, A2 => n19606, B1 => n19619, B2 => 
                           n2359, ZN => n7486);
   U6408 : OAI22_X1 port map( A1 => n20403, A2 => n19605, B1 => n19618, B2 => 
                           n2358, ZN => n7487);
   U6409 : OAI22_X1 port map( A1 => n20406, A2 => n19605, B1 => n19618, B2 => 
                           n2357, ZN => n7488);
   U6410 : OAI22_X1 port map( A1 => n20409, A2 => n19605, B1 => n19618, B2 => 
                           n2356, ZN => n7489);
   U6411 : OAI22_X1 port map( A1 => n20412, A2 => n19605, B1 => n19618, B2 => 
                           n2355, ZN => n7490);
   U6412 : OAI22_X1 port map( A1 => n20415, A2 => n19605, B1 => n19617, B2 => 
                           n2354, ZN => n7491);
   U6413 : OAI22_X1 port map( A1 => n20418, A2 => n19605, B1 => n19617, B2 => 
                           n2353, ZN => n7492);
   U6414 : OAI22_X1 port map( A1 => n20421, A2 => n19605, B1 => n19617, B2 => 
                           n2352, ZN => n7493);
   U6415 : OAI22_X1 port map( A1 => n20424, A2 => n19605, B1 => n19617, B2 => 
                           n2351, ZN => n7494);
   U6416 : OAI22_X1 port map( A1 => n20427, A2 => n19605, B1 => n19616, B2 => 
                           n2350, ZN => n7495);
   U6417 : OAI22_X1 port map( A1 => n20430, A2 => n19605, B1 => n19616, B2 => 
                           n2349, ZN => n7496);
   U6418 : OAI22_X1 port map( A1 => n20433, A2 => n19605, B1 => n19616, B2 => 
                           n2348, ZN => n7497);
   U6419 : OAI22_X1 port map( A1 => n20436, A2 => n19605, B1 => n19616, B2 => 
                           n2347, ZN => n7498);
   U6420 : OAI22_X1 port map( A1 => n20439, A2 => n19604, B1 => n19615, B2 => 
                           n2346, ZN => n7499);
   U6421 : OAI22_X1 port map( A1 => n20442, A2 => n19604, B1 => n19615, B2 => 
                           n2345, ZN => n7500);
   U6422 : OAI22_X1 port map( A1 => n20445, A2 => n19604, B1 => n19615, B2 => 
                           n2344, ZN => n7501);
   U6423 : OAI22_X1 port map( A1 => n20448, A2 => n19604, B1 => n19615, B2 => 
                           n2343, ZN => n7502);
   U6424 : OAI22_X1 port map( A1 => n20451, A2 => n19604, B1 => n19614, B2 => 
                           n2342, ZN => n7503);
   U6425 : OAI22_X1 port map( A1 => n20454, A2 => n19604, B1 => n19614, B2 => 
                           n2341, ZN => n7504);
   U6426 : OAI22_X1 port map( A1 => n20457, A2 => n19604, B1 => n19614, B2 => 
                           n2340, ZN => n7505);
   U6427 : OAI22_X1 port map( A1 => n20460, A2 => n19604, B1 => n19614, B2 => 
                           n2339, ZN => n7506);
   U6428 : OAI22_X1 port map( A1 => n20463, A2 => n19604, B1 => n19613, B2 => 
                           n2338, ZN => n7507);
   U6429 : OAI22_X1 port map( A1 => n20466, A2 => n19604, B1 => n19613, B2 => 
                           n2337, ZN => n7508);
   U6430 : OAI22_X1 port map( A1 => n20469, A2 => n19604, B1 => n19613, B2 => 
                           n2336, ZN => n7509);
   U6431 : OAI22_X1 port map( A1 => n20472, A2 => n19604, B1 => n19613, B2 => 
                           n2333, ZN => n7510);
   U6432 : OAI22_X1 port map( A1 => n20475, A2 => n19606, B1 => n19612, B2 => 
                           n2330, ZN => n7511);
   U6433 : OAI22_X1 port map( A1 => n20478, A2 => n19605, B1 => n19612, B2 => 
                           n2327, ZN => n7512);
   U6434 : OAI22_X1 port map( A1 => n20481, A2 => n19604, B1 => n19612, B2 => 
                           n2324, ZN => n7513);
   U6435 : OAI22_X1 port map( A1 => n20484, A2 => n19606, B1 => n19612, B2 => 
                           n2321, ZN => n7514);
   U6436 : OAI22_X1 port map( A1 => n20487, A2 => n19605, B1 => n19611, B2 => 
                           n2318, ZN => n7515);
   U6437 : OAI22_X1 port map( A1 => n20490, A2 => n19604, B1 => n19611, B2 => 
                           n2315, ZN => n7516);
   U6438 : OAI22_X1 port map( A1 => n20493, A2 => n19606, B1 => n19611, B2 => 
                           n2312, ZN => n7517);
   U6439 : OAI22_X1 port map( A1 => n20496, A2 => n19605, B1 => n19611, B2 => 
                           n2309, ZN => n7518);
   U6440 : OAI22_X1 port map( A1 => n20499, A2 => n19604, B1 => n19610, B2 => 
                           n2306, ZN => n7519);
   U6441 : OAI22_X1 port map( A1 => n20502, A2 => n19606, B1 => n19610, B2 => 
                           n2303, ZN => n7520);
   U6442 : OAI22_X1 port map( A1 => n20505, A2 => n19605, B1 => n19610, B2 => 
                           n2300, ZN => n7521);
   U6443 : OAI22_X1 port map( A1 => n20508, A2 => n19605, B1 => n19610, B2 => 
                           n2297, ZN => n7522);
   U6444 : OAI22_X1 port map( A1 => n20511, A2 => n19606, B1 => n19609, B2 => 
                           n2294, ZN => n7523);
   U6445 : OAI22_X1 port map( A1 => n20514, A2 => n19605, B1 => n19609, B2 => 
                           n2291, ZN => n7524);
   U6446 : OAI22_X1 port map( A1 => n20517, A2 => n19604, B1 => n19609, B2 => 
                           n2288, ZN => n7525);
   U6447 : OAI22_X1 port map( A1 => n20520, A2 => n19604, B1 => n19609, B2 => 
                           n2285, ZN => n7526);
   U6448 : OAI22_X1 port map( A1 => n20523, A2 => n19606, B1 => n19608, B2 => 
                           n2282, ZN => n7527);
   U6449 : OAI22_X1 port map( A1 => n20526, A2 => n19605, B1 => n19608, B2 => 
                           n2279, ZN => n7528);
   U6450 : OAI22_X1 port map( A1 => n20529, A2 => n19604, B1 => n19608, B2 => 
                           n2276, ZN => n7529);
   U6451 : OAI22_X1 port map( A1 => n20532, A2 => n19606, B1 => n19608, B2 => 
                           n2273, ZN => n7530);
   U6452 : OAI22_X1 port map( A1 => n20535, A2 => n19606, B1 => n19607, B2 => 
                           n2270, ZN => n7531);
   U6453 : OAI22_X1 port map( A1 => n20538, A2 => n19605, B1 => n19607, B2 => 
                           n2267, ZN => n7532);
   U6454 : OAI22_X1 port map( A1 => n20541, A2 => n19604, B1 => n19607, B2 => 
                           n2264, ZN => n7533);
   U6455 : OAI22_X1 port map( A1 => n20572, A2 => n19605, B1 => n19607, B2 => 
                           n2261, ZN => n7534);
   U6456 : OAI22_X1 port map( A1 => n20356, A2 => n19913, B1 => n19930, B2 => 
                           n2013, ZN => n8175);
   U6457 : OAI22_X1 port map( A1 => n20359, A2 => n19912, B1 => n19930, B2 => 
                           n2012, ZN => n8176);
   U6458 : OAI22_X1 port map( A1 => n20362, A2 => n19912, B1 => n19930, B2 => 
                           n2011, ZN => n8177);
   U6459 : OAI22_X1 port map( A1 => n20365, A2 => n19914, B1 => n19930, B2 => 
                           n2010, ZN => n8178);
   U6460 : OAI22_X1 port map( A1 => n20355, A2 => n19605, B1 => n19622, B2 => 
                           n2374, ZN => n7471);
   U6461 : OAI22_X1 port map( A1 => n20358, A2 => n19604, B1 => n19622, B2 => 
                           n2373, ZN => n7472);
   U6462 : OAI22_X1 port map( A1 => n20361, A2 => n19604, B1 => n19622, B2 => 
                           n2372, ZN => n7473);
   U6463 : OAI22_X1 port map( A1 => n20364, A2 => n19606, B1 => n19622, B2 => 
                           n2371, ZN => n7474);
   U6464 : OAI22_X1 port map( A1 => n20368, A2 => n19886, B1 => n19901, B2 => 
                           n2077, ZN => n8115);
   U6465 : OAI22_X1 port map( A1 => n20371, A2 => n19886, B1 => n19901, B2 => 
                           n2076, ZN => n8116);
   U6466 : OAI22_X1 port map( A1 => n20374, A2 => n19886, B1 => n19901, B2 => 
                           n2075, ZN => n8117);
   U6467 : OAI22_X1 port map( A1 => n20377, A2 => n19886, B1 => n19901, B2 => 
                           n2074, ZN => n8118);
   U6468 : OAI22_X1 port map( A1 => n20380, A2 => n19886, B1 => n19900, B2 => 
                           n2073, ZN => n8119);
   U6469 : OAI22_X1 port map( A1 => n20383, A2 => n19886, B1 => n19900, B2 => 
                           n2072, ZN => n8120);
   U6470 : OAI22_X1 port map( A1 => n20386, A2 => n19886, B1 => n19900, B2 => 
                           n2071, ZN => n8121);
   U6471 : OAI22_X1 port map( A1 => n20389, A2 => n19886, B1 => n19900, B2 => 
                           n2070, ZN => n8122);
   U6472 : OAI22_X1 port map( A1 => n20392, A2 => n19886, B1 => n19899, B2 => 
                           n2069, ZN => n8123);
   U6473 : OAI22_X1 port map( A1 => n20395, A2 => n19886, B1 => n19899, B2 => 
                           n2068, ZN => n8124);
   U6474 : OAI22_X1 port map( A1 => n20398, A2 => n19886, B1 => n19899, B2 => 
                           n2067, ZN => n8125);
   U6475 : OAI22_X1 port map( A1 => n20401, A2 => n19886, B1 => n19899, B2 => 
                           n2066, ZN => n8126);
   U6476 : OAI22_X1 port map( A1 => n20404, A2 => n19885, B1 => n19898, B2 => 
                           n2065, ZN => n8127);
   U6477 : OAI22_X1 port map( A1 => n20407, A2 => n19885, B1 => n19898, B2 => 
                           n2064, ZN => n8128);
   U6478 : OAI22_X1 port map( A1 => n20410, A2 => n19885, B1 => n19898, B2 => 
                           n2063, ZN => n8129);
   U6479 : OAI22_X1 port map( A1 => n20413, A2 => n19885, B1 => n19898, B2 => 
                           n2062, ZN => n8130);
   U6480 : OAI22_X1 port map( A1 => n20416, A2 => n19885, B1 => n19897, B2 => 
                           n2061, ZN => n8131);
   U6481 : OAI22_X1 port map( A1 => n20419, A2 => n19885, B1 => n19897, B2 => 
                           n2060, ZN => n8132);
   U6482 : OAI22_X1 port map( A1 => n20422, A2 => n19885, B1 => n19897, B2 => 
                           n2059, ZN => n8133);
   U6483 : OAI22_X1 port map( A1 => n20425, A2 => n19885, B1 => n19897, B2 => 
                           n2058, ZN => n8134);
   U6484 : OAI22_X1 port map( A1 => n20428, A2 => n19885, B1 => n19896, B2 => 
                           n2057, ZN => n8135);
   U6485 : OAI22_X1 port map( A1 => n20431, A2 => n19885, B1 => n19896, B2 => 
                           n2056, ZN => n8136);
   U6486 : OAI22_X1 port map( A1 => n20434, A2 => n19885, B1 => n19896, B2 => 
                           n2055, ZN => n8137);
   U6487 : OAI22_X1 port map( A1 => n20437, A2 => n19885, B1 => n19896, B2 => 
                           n2054, ZN => n8138);
   U6488 : OAI22_X1 port map( A1 => n20440, A2 => n19884, B1 => n19895, B2 => 
                           n2053, ZN => n8139);
   U6489 : OAI22_X1 port map( A1 => n20443, A2 => n19884, B1 => n19895, B2 => 
                           n2052, ZN => n8140);
   U6490 : OAI22_X1 port map( A1 => n20446, A2 => n19884, B1 => n19895, B2 => 
                           n2051, ZN => n8141);
   U6491 : OAI22_X1 port map( A1 => n20449, A2 => n19884, B1 => n19895, B2 => 
                           n2050, ZN => n8142);
   U6492 : OAI22_X1 port map( A1 => n20452, A2 => n19884, B1 => n19894, B2 => 
                           n2049, ZN => n8143);
   U6493 : OAI22_X1 port map( A1 => n20455, A2 => n19884, B1 => n19894, B2 => 
                           n2048, ZN => n8144);
   U6494 : OAI22_X1 port map( A1 => n20458, A2 => n19884, B1 => n19894, B2 => 
                           n2047, ZN => n8145);
   U6495 : OAI22_X1 port map( A1 => n20461, A2 => n19884, B1 => n19894, B2 => 
                           n2046, ZN => n8146);
   U6496 : OAI22_X1 port map( A1 => n20464, A2 => n19884, B1 => n19893, B2 => 
                           n2045, ZN => n8147);
   U6497 : OAI22_X1 port map( A1 => n20467, A2 => n19884, B1 => n19893, B2 => 
                           n2044, ZN => n8148);
   U6498 : OAI22_X1 port map( A1 => n20470, A2 => n19884, B1 => n19893, B2 => 
                           n2043, ZN => n8149);
   U6499 : OAI22_X1 port map( A1 => n20473, A2 => n19884, B1 => n19893, B2 => 
                           n2042, ZN => n8150);
   U6500 : OAI22_X1 port map( A1 => n20476, A2 => n19886, B1 => n19892, B2 => 
                           n2041, ZN => n8151);
   U6501 : OAI22_X1 port map( A1 => n20479, A2 => n19885, B1 => n19892, B2 => 
                           n2040, ZN => n8152);
   U6502 : OAI22_X1 port map( A1 => n20482, A2 => n19884, B1 => n19892, B2 => 
                           n2039, ZN => n8153);
   U6503 : OAI22_X1 port map( A1 => n20485, A2 => n19886, B1 => n19892, B2 => 
                           n2038, ZN => n8154);
   U6504 : OAI22_X1 port map( A1 => n20488, A2 => n19885, B1 => n19891, B2 => 
                           n2037, ZN => n8155);
   U6505 : OAI22_X1 port map( A1 => n20491, A2 => n19884, B1 => n19891, B2 => 
                           n2036, ZN => n8156);
   U6506 : OAI22_X1 port map( A1 => n20494, A2 => n19886, B1 => n19891, B2 => 
                           n2035, ZN => n8157);
   U6507 : OAI22_X1 port map( A1 => n20497, A2 => n19885, B1 => n19891, B2 => 
                           n2034, ZN => n8158);
   U6508 : OAI22_X1 port map( A1 => n20500, A2 => n19884, B1 => n19890, B2 => 
                           n2033, ZN => n8159);
   U6509 : OAI22_X1 port map( A1 => n20503, A2 => n19886, B1 => n19890, B2 => 
                           n2032, ZN => n8160);
   U6510 : OAI22_X1 port map( A1 => n20506, A2 => n19885, B1 => n19890, B2 => 
                           n2031, ZN => n8161);
   U6511 : OAI22_X1 port map( A1 => n20509, A2 => n19885, B1 => n19890, B2 => 
                           n2030, ZN => n8162);
   U6512 : OAI22_X1 port map( A1 => n20512, A2 => n19886, B1 => n19889, B2 => 
                           n2029, ZN => n8163);
   U6513 : OAI22_X1 port map( A1 => n20515, A2 => n19885, B1 => n19889, B2 => 
                           n2028, ZN => n8164);
   U6514 : OAI22_X1 port map( A1 => n20518, A2 => n19884, B1 => n19889, B2 => 
                           n2027, ZN => n8165);
   U6515 : OAI22_X1 port map( A1 => n20521, A2 => n19884, B1 => n19889, B2 => 
                           n2026, ZN => n8166);
   U6516 : OAI22_X1 port map( A1 => n20524, A2 => n19886, B1 => n19888, B2 => 
                           n2025, ZN => n8167);
   U6517 : OAI22_X1 port map( A1 => n20527, A2 => n19885, B1 => n19888, B2 => 
                           n2024, ZN => n8168);
   U6518 : OAI22_X1 port map( A1 => n20530, A2 => n19884, B1 => n19888, B2 => 
                           n2023, ZN => n8169);
   U6519 : OAI22_X1 port map( A1 => n20533, A2 => n19886, B1 => n19888, B2 => 
                           n2022, ZN => n8170);
   U6520 : OAI22_X1 port map( A1 => n20536, A2 => n19886, B1 => n19887, B2 => 
                           n2021, ZN => n8171);
   U6521 : OAI22_X1 port map( A1 => n20539, A2 => n19885, B1 => n19887, B2 => 
                           n2020, ZN => n8172);
   U6522 : OAI22_X1 port map( A1 => n20542, A2 => n19884, B1 => n19887, B2 => 
                           n2019, ZN => n8173);
   U6523 : OAI22_X1 port map( A1 => n20573, A2 => n19885, B1 => n19887, B2 => 
                           n2018, ZN => n8174);
   U6524 : OAI22_X1 port map( A1 => n20356, A2 => n19885, B1 => n19902, B2 => 
                           n2081, ZN => n8111);
   U6525 : OAI22_X1 port map( A1 => n20359, A2 => n19884, B1 => n19902, B2 => 
                           n2080, ZN => n8112);
   U6526 : OAI22_X1 port map( A1 => n20362, A2 => n19884, B1 => n19902, B2 => 
                           n2079, ZN => n8113);
   U6527 : OAI22_X1 port map( A1 => n20365, A2 => n19886, B1 => n19902, B2 => 
                           n2078, ZN => n8114);
   U6528 : NAND4_X1 port map( A1 => n11559, A2 => n11560, A3 => rd1, A4 => 
                           n11561, ZN => n2222);
   U6529 : NAND2_X1 port map( A1 => N150, A2 => n11565, ZN => n11560);
   U6530 : AOI221_X1 port map( B1 => n2228, B2 => n11562, C1 => n1940, C2 => 
                           n11563, A => n11564, ZN => n11561);
   U6531 : OAI22_X1 port map( A1 => N79, A2 => n1947, B1 => N78, B2 => n2094, 
                           ZN => n11564);
   U6532 : NAND4_X1 port map( A1 => n5321, A2 => n5322, A3 => n5323, A4 => 
                           n5324, ZN => n7263);
   U6533 : AOI222_X1 port map( A1 => out_to_mem_60_port, A2 => n18917, B1 => 
                           n18914, B2 => n18176, C1 => registers_3_60_port, C2 
                           => n18908, ZN => n5321);
   U6534 : AOI221_X1 port map( B1 => n18941, B2 => n5337, C1 => n18935, C2 => 
                           n5338, A => n5339, ZN => n5322);
   U6535 : AOI211_X1 port map( C1 => registers_4_60_port, C2 => n18983, A => 
                           n5333, B => n5334, ZN => n5323);
   U6536 : NAND4_X1 port map( A1 => n4516, A2 => n4581, A3 => n4582, A4 => 
                           n4583, ZN => n7267);
   U6537 : AOI222_X1 port map( A1 => out_to_mem_61_port, A2 => n18917, B1 => 
                           n18914, B2 => n18177, C1 => registers_3_61_port, C2 
                           => n18908, ZN => n4516);
   U6538 : AOI221_X1 port map( B1 => n18941, B2 => n4852, C1 => n18935, C2 => 
                           n4853, A => n4854, ZN => n4581);
   U6539 : AOI211_X1 port map( C1 => registers_4_61_port, C2 => n18983, A => 
                           n4784, B => n4785, ZN => n4582);
   U6540 : NAND4_X1 port map( A1 => n3298, A2 => n3299, A3 => n3300, A4 => 
                           n3301, ZN => n7271);
   U6541 : AOI222_X1 port map( A1 => out_to_mem_62_port, A2 => n18917, B1 => 
                           n18914, B2 => n18178, C1 => registers_3_62_port, C2 
                           => n18908, ZN => n3298);
   U6542 : AOI221_X1 port map( B1 => n18941, B2 => n3570, C1 => n18935, C2 => 
                           n3571, A => n3572, ZN => n3299);
   U6543 : AOI211_X1 port map( C1 => registers_4_62_port, C2 => n18983, A => 
                           n3438, B => n3503, ZN => n3300);
   U6544 : NAND4_X1 port map( A1 => n3139, A2 => n3140, A3 => n3141, A4 => 
                           n3142, ZN => n7275);
   U6545 : AOI222_X1 port map( A1 => out_to_mem_63_port, A2 => n18916, B1 => 
                           n18914, B2 => n18179, C1 => registers_3_63_port, C2 
                           => n18908, ZN => n3139);
   U6546 : AOI221_X1 port map( B1 => n18941, B2 => n3188, C1 => n18935, C2 => 
                           n3192, A => n3194, ZN => n3140);
   U6547 : AOI211_X1 port map( C1 => registers_4_63_port, C2 => n18983, A => 
                           n3167, B => n3168, ZN => n3141);
   U6548 : NAND4_X1 port map( A1 => n6807, A2 => n6808, A3 => n6809, A4 => 
                           n6810, ZN => n7175);
   U6549 : AOI222_X1 port map( A1 => out_to_mem_38_port, A2 => n18915, B1 => 
                           n18912, B2 => n18180, C1 => registers_3_38_port, C2 
                           => n18906, ZN => n6807);
   U6550 : AOI221_X1 port map( B1 => n18939, B2 => n6823, C1 => n18933, C2 => 
                           n6824, A => n6825, ZN => n6808);
   U6551 : NAND4_X1 port map( A1 => n6739, A2 => n6740, A3 => n6741, A4 => 
                           n6742, ZN => n7179);
   U6552 : AOI222_X1 port map( A1 => out_to_mem_39_port, A2 => n18915, B1 => 
                           n18912, B2 => n18181, C1 => registers_3_39_port, C2 
                           => n18906, ZN => n6739);
   U6553 : AOI221_X1 port map( B1 => n18939, B2 => n6756, C1 => n18933, C2 => 
                           n6757, A => n6758, ZN => n6740);
   U6554 : AOI211_X1 port map( C1 => registers_4_39_port, C2 => n18981, A => 
                           n6752, B => n6753, ZN => n6741);
   U6555 : NAND4_X1 port map( A1 => n6672, A2 => n6673, A3 => n6674, A4 => 
                           n6675, ZN => n7183);
   U6556 : AOI222_X1 port map( A1 => out_to_mem_40_port, A2 => n18915, B1 => 
                           n18912, B2 => n18182, C1 => registers_3_40_port, C2 
                           => n18906, ZN => n6672);
   U6557 : AOI221_X1 port map( B1 => n18939, B2 => n6688, C1 => n18933, C2 => 
                           n6689, A => n6690, ZN => n6673);
   U6558 : AOI211_X1 port map( C1 => registers_4_40_port, C2 => n18981, A => 
                           n6684, B => n6685, ZN => n6674);
   U6559 : NAND4_X1 port map( A1 => n6605, A2 => n6606, A3 => n6607, A4 => 
                           n6608, ZN => n7187);
   U6560 : AOI222_X1 port map( A1 => out_to_mem_41_port, A2 => n18915, B1 => 
                           n18912, B2 => n18183, C1 => registers_3_41_port, C2 
                           => n18906, ZN => n6605);
   U6561 : AOI221_X1 port map( B1 => n18939, B2 => n6621, C1 => n18933, C2 => 
                           n6622, A => n6623, ZN => n6606);
   U6562 : AOI211_X1 port map( C1 => registers_4_41_port, C2 => n18981, A => 
                           n6617, B => n6618, ZN => n6607);
   U6563 : NAND4_X1 port map( A1 => n6539, A2 => n6540, A3 => n6541, A4 => 
                           n6542, ZN => n7191);
   U6564 : AOI222_X1 port map( A1 => out_to_mem_42_port, A2 => n18915, B1 => 
                           n18912, B2 => n18184, C1 => registers_3_42_port, C2 
                           => n18906, ZN => n6539);
   U6565 : AOI221_X1 port map( B1 => n18939, B2 => n6555, C1 => n18933, C2 => 
                           n6556, A => n6557, ZN => n6540);
   U6566 : AOI211_X1 port map( C1 => registers_4_42_port, C2 => n18981, A => 
                           n6551, B => n6552, ZN => n6541);
   U6567 : NAND4_X1 port map( A1 => n6473, A2 => n6474, A3 => n6475, A4 => 
                           n6476, ZN => n7195);
   U6568 : AOI222_X1 port map( A1 => out_to_mem_43_port, A2 => n18915, B1 => 
                           n18912, B2 => n18185, C1 => registers_3_43_port, C2 
                           => n18906, ZN => n6473);
   U6569 : AOI221_X1 port map( B1 => n18939, B2 => n6489, C1 => n18933, C2 => 
                           n6490, A => n6491, ZN => n6474);
   U6570 : AOI211_X1 port map( C1 => registers_4_43_port, C2 => n18981, A => 
                           n6485, B => n6486, ZN => n6475);
   U6571 : NAND4_X1 port map( A1 => n6407, A2 => n6408, A3 => n6409, A4 => 
                           n6410, ZN => n7199);
   U6572 : AOI222_X1 port map( A1 => out_to_mem_44_port, A2 => n18915, B1 => 
                           n18912, B2 => n18186, C1 => registers_3_44_port, C2 
                           => n18906, ZN => n6407);
   U6573 : AOI221_X1 port map( B1 => n18939, B2 => n6423, C1 => n18933, C2 => 
                           n6424, A => n6425, ZN => n6408);
   U6574 : AOI211_X1 port map( C1 => registers_4_44_port, C2 => n18981, A => 
                           n6419, B => n6420, ZN => n6409);
   U6575 : NAND4_X1 port map( A1 => n6341, A2 => n6342, A3 => n6343, A4 => 
                           n6344, ZN => n7203);
   U6576 : AOI222_X1 port map( A1 => out_to_mem_45_port, A2 => n18915, B1 => 
                           n18912, B2 => n18187, C1 => registers_3_45_port, C2 
                           => n18906, ZN => n6341);
   U6577 : AOI221_X1 port map( B1 => n18939, B2 => n6357, C1 => n18933, C2 => 
                           n6358, A => n6359, ZN => n6342);
   U6578 : AOI211_X1 port map( C1 => registers_4_45_port, C2 => n18981, A => 
                           n6353, B => n6354, ZN => n6343);
   U6579 : NAND4_X1 port map( A1 => n6275, A2 => n6276, A3 => n6277, A4 => 
                           n6278, ZN => n7207);
   U6580 : AOI222_X1 port map( A1 => out_to_mem_46_port, A2 => n18915, B1 => 
                           n18912, B2 => n18188, C1 => registers_3_46_port, C2 
                           => n18906, ZN => n6275);
   U6581 : AOI221_X1 port map( B1 => n18939, B2 => n6291, C1 => n18933, C2 => 
                           n6292, A => n6293, ZN => n6276);
   U6582 : AOI211_X1 port map( C1 => registers_4_46_port, C2 => n18981, A => 
                           n6287, B => n6288, ZN => n6277);
   U6583 : NAND4_X1 port map( A1 => n6209, A2 => n6210, A3 => n6211, A4 => 
                           n6212, ZN => n7211);
   U6584 : AOI222_X1 port map( A1 => out_to_mem_47_port, A2 => n18915, B1 => 
                           n18912, B2 => n18189, C1 => registers_3_47_port, C2 
                           => n18906, ZN => n6209);
   U6585 : AOI221_X1 port map( B1 => n18939, B2 => n6225, C1 => n18933, C2 => 
                           n6226, A => n6227, ZN => n6210);
   U6586 : AOI211_X1 port map( C1 => registers_4_47_port, C2 => n18981, A => 
                           n6221, B => n6222, ZN => n6211);
   U6587 : NAND4_X1 port map( A1 => n6143, A2 => n6144, A3 => n6145, A4 => 
                           n6146, ZN => n7215);
   U6588 : AOI222_X1 port map( A1 => out_to_mem_48_port, A2 => n18915, B1 => 
                           n18913, B2 => n18190, C1 => registers_3_48_port, C2 
                           => n18907, ZN => n6143);
   U6589 : AOI221_X1 port map( B1 => n18940, B2 => n6159, C1 => n18934, C2 => 
                           n6160, A => n6161, ZN => n6144);
   U6590 : AOI211_X1 port map( C1 => registers_4_48_port, C2 => n18982, A => 
                           n6155, B => n6156, ZN => n6145);
   U6591 : NAND4_X1 port map( A1 => n6077, A2 => n6078, A3 => n6079, A4 => 
                           n6080, ZN => n7219);
   U6592 : AOI222_X1 port map( A1 => out_to_mem_49_port, A2 => n18915, B1 => 
                           n18913, B2 => n18191, C1 => registers_3_49_port, C2 
                           => n18907, ZN => n6077);
   U6593 : AOI221_X1 port map( B1 => n18940, B2 => n6093, C1 => n18934, C2 => 
                           n6094, A => n6095, ZN => n6078);
   U6594 : AOI211_X1 port map( C1 => registers_4_49_port, C2 => n18982, A => 
                           n6089, B => n6090, ZN => n6079);
   U6595 : NAND4_X1 port map( A1 => n6009, A2 => n6010, A3 => n6011, A4 => 
                           n6012, ZN => n7223);
   U6596 : AOI222_X1 port map( A1 => out_to_mem_50_port, A2 => n18915, B1 => 
                           n18913, B2 => n18192, C1 => registers_3_50_port, C2 
                           => n18907, ZN => n6009);
   U6597 : AOI221_X1 port map( B1 => n18940, B2 => n6025, C1 => n18934, C2 => 
                           n6026, A => n6027, ZN => n6010);
   U6598 : AOI211_X1 port map( C1 => registers_4_50_port, C2 => n18982, A => 
                           n6021, B => n6022, ZN => n6011);
   U6599 : NAND4_X1 port map( A1 => n5941, A2 => n5942, A3 => n5943, A4 => 
                           n5944, ZN => n7227);
   U6600 : AOI222_X1 port map( A1 => out_to_mem_51_port, A2 => n18915, B1 => 
                           n18913, B2 => n18193, C1 => registers_3_51_port, C2 
                           => n18907, ZN => n5941);
   U6601 : AOI221_X1 port map( B1 => n18940, B2 => n5957, C1 => n18934, C2 => 
                           n5958, A => n5959, ZN => n5942);
   U6602 : AOI211_X1 port map( C1 => registers_4_51_port, C2 => n18982, A => 
                           n5953, B => n5954, ZN => n5943);
   U6603 : NAND4_X1 port map( A1 => n5874, A2 => n5875, A3 => n5876, A4 => 
                           n5877, ZN => n7231);
   U6604 : AOI222_X1 port map( A1 => out_to_mem_52_port, A2 => n18915, B1 => 
                           n18913, B2 => n18194, C1 => registers_3_52_port, C2 
                           => n18907, ZN => n5874);
   U6605 : AOI221_X1 port map( B1 => n18940, B2 => n5890, C1 => n18934, C2 => 
                           n5891, A => n5892, ZN => n5875);
   U6606 : AOI211_X1 port map( C1 => registers_4_52_port, C2 => n18982, A => 
                           n5886, B => n5887, ZN => n5876);
   U6607 : NAND4_X1 port map( A1 => n5807, A2 => n5808, A3 => n5809, A4 => 
                           n5810, ZN => n7235);
   U6608 : AOI222_X1 port map( A1 => out_to_mem_53_port, A2 => n18915, B1 => 
                           n18913, B2 => n18195, C1 => registers_3_53_port, C2 
                           => n18907, ZN => n5807);
   U6609 : AOI221_X1 port map( B1 => n18940, B2 => n5823, C1 => n18934, C2 => 
                           n5824, A => n5825, ZN => n5808);
   U6610 : AOI211_X1 port map( C1 => registers_4_53_port, C2 => n18982, A => 
                           n5819, B => n5820, ZN => n5809);
   U6611 : NAND4_X1 port map( A1 => n5735, A2 => n5736, A3 => n5737, A4 => 
                           n5738, ZN => n7239);
   U6612 : AOI222_X1 port map( A1 => out_to_mem_54_port, A2 => n18915, B1 => 
                           n18913, B2 => n18196, C1 => registers_3_54_port, C2 
                           => n18907, ZN => n5735);
   U6613 : AOI221_X1 port map( B1 => n18940, B2 => n5751, C1 => n18934, C2 => 
                           n5752, A => n5753, ZN => n5736);
   U6614 : AOI211_X1 port map( C1 => registers_4_54_port, C2 => n18982, A => 
                           n5747, B => n5748, ZN => n5737);
   U6615 : NAND4_X1 port map( A1 => n5665, A2 => n5666, A3 => n5667, A4 => 
                           n5668, ZN => n7243);
   U6616 : AOI222_X1 port map( A1 => out_to_mem_55_port, A2 => n18915, B1 => 
                           n18913, B2 => n18197, C1 => registers_3_55_port, C2 
                           => n18907, ZN => n5665);
   U6617 : AOI221_X1 port map( B1 => n18940, B2 => n5681, C1 => n18934, C2 => 
                           n5682, A => n5683, ZN => n5666);
   U6618 : AOI211_X1 port map( C1 => registers_4_55_port, C2 => n18982, A => 
                           n5677, B => n5678, ZN => n5667);
   U6619 : NAND4_X1 port map( A1 => n5597, A2 => n5598, A3 => n5599, A4 => 
                           n5600, ZN => n7247);
   U6620 : AOI222_X1 port map( A1 => out_to_mem_56_port, A2 => n18915, B1 => 
                           n18913, B2 => n18198, C1 => registers_3_56_port, C2 
                           => n18907, ZN => n5597);
   U6621 : AOI221_X1 port map( B1 => n18940, B2 => n5613, C1 => n18934, C2 => 
                           n5614, A => n5615, ZN => n5598);
   U6622 : AOI211_X1 port map( C1 => registers_4_56_port, C2 => n18982, A => 
                           n5609, B => n5610, ZN => n5599);
   U6623 : NAND4_X1 port map( A1 => n5528, A2 => n5529, A3 => n5530, A4 => 
                           n5531, ZN => n7251);
   U6624 : AOI222_X1 port map( A1 => out_to_mem_57_port, A2 => n18917, B1 => 
                           n18913, B2 => n18199, C1 => registers_3_57_port, C2 
                           => n18907, ZN => n5528);
   U6625 : AOI221_X1 port map( B1 => n18940, B2 => n5544, C1 => n18934, C2 => 
                           n5545, A => n5546, ZN => n5529);
   U6626 : AOI211_X1 port map( C1 => registers_4_57_port, C2 => n18982, A => 
                           n5540, B => n5541, ZN => n5530);
   U6627 : NAND4_X1 port map( A1 => n5459, A2 => n5460, A3 => n5461, A4 => 
                           n5462, ZN => n7255);
   U6628 : AOI222_X1 port map( A1 => out_to_mem_58_port, A2 => n18917, B1 => 
                           n18913, B2 => n18200, C1 => registers_3_58_port, C2 
                           => n18907, ZN => n5459);
   U6629 : AOI221_X1 port map( B1 => n18940, B2 => n5475, C1 => n18934, C2 => 
                           n5476, A => n5477, ZN => n5460);
   U6630 : AOI211_X1 port map( C1 => registers_4_58_port, C2 => n18982, A => 
                           n5471, B => n5472, ZN => n5461);
   U6631 : NAND4_X1 port map( A1 => n5391, A2 => n5392, A3 => n5393, A4 => 
                           n5394, ZN => n7259);
   U6632 : AOI222_X1 port map( A1 => out_to_mem_59_port, A2 => n18917, B1 => 
                           n18913, B2 => n18201, C1 => registers_3_59_port, C2 
                           => n18907, ZN => n5391);
   U6633 : AOI221_X1 port map( B1 => n18940, B2 => n5407, C1 => n18934, C2 => 
                           n5408, A => n5409, ZN => n5392);
   U6634 : AOI211_X1 port map( C1 => registers_4_59_port, C2 => n18982, A => 
                           n5403, B => n5404, ZN => n5393);
   U6635 : NAND4_X1 port map( A1 => n11662, A2 => n11663, A3 => n11664, A4 => 
                           n11665, ZN => n7023);
   U6636 : AOI222_X1 port map( A1 => out_to_mem_0_port, A2 => n18917, B1 => 
                           n18909, B2 => n11719, C1 => registers_3_0_port, C2 
                           => n18903, ZN => n11662);
   U6637 : AOI221_X1 port map( B1 => n18936, B2 => n11712, C1 => n18930, C2 => 
                           n11713, A => n11714, ZN => n11663);
   U6638 : AOI211_X1 port map( C1 => registers_4_0_port, C2 => n18978, A => 
                           n11697, B => n11698, ZN => n11664);
   U6639 : NAND4_X1 port map( A1 => n11534, A2 => n11535, A3 => n11536, A4 => 
                           n11537, ZN => n7027);
   U6640 : AOI222_X1 port map( A1 => out_to_mem_1_port, A2 => n18916, B1 => 
                           n18909, B2 => n11554, C1 => registers_3_1_port, C2 
                           => n18903, ZN => n11534);
   U6641 : AOI221_X1 port map( B1 => n18936, B2 => n11551, C1 => n18930, C2 => 
                           n11552, A => n11553, ZN => n11535);
   U6642 : AOI211_X1 port map( C1 => registers_4_1_port, C2 => n18978, A => 
                           n11547, B => n11548, ZN => n11536);
   U6643 : NAND4_X1 port map( A1 => n11467, A2 => n11468, A3 => n11469, A4 => 
                           n11470, ZN => n7031);
   U6644 : AOI222_X1 port map( A1 => out_to_mem_2_port, A2 => n18916, B1 => 
                           n18909, B2 => n11486, C1 => registers_3_2_port, C2 
                           => n18903, ZN => n11467);
   U6645 : AOI221_X1 port map( B1 => n18936, B2 => n11483, C1 => n18930, C2 => 
                           n11484, A => n11485, ZN => n11468);
   U6646 : AOI211_X1 port map( C1 => registers_4_2_port, C2 => n18978, A => 
                           n11479, B => n11480, ZN => n11469);
   U6647 : NAND4_X1 port map( A1 => n11400, A2 => n11401, A3 => n11402, A4 => 
                           n11403, ZN => n7035);
   U6648 : AOI222_X1 port map( A1 => out_to_mem_3_port, A2 => n18915, B1 => 
                           n18909, B2 => n11419, C1 => registers_3_3_port, C2 
                           => n18903, ZN => n11400);
   U6649 : AOI221_X1 port map( B1 => n18936, B2 => n11416, C1 => n18930, C2 => 
                           n11417, A => n11418, ZN => n11401);
   U6650 : AOI211_X1 port map( C1 => registers_4_3_port, C2 => n18978, A => 
                           n11412, B => n11413, ZN => n11402);
   U6651 : NAND4_X1 port map( A1 => n11333, A2 => n11334, A3 => n11335, A4 => 
                           n11336, ZN => n7039);
   U6652 : AOI222_X1 port map( A1 => out_to_mem_4_port, A2 => n18917, B1 => 
                           n18909, B2 => n18202, C1 => registers_3_4_port, C2 
                           => n18903, ZN => n11333);
   U6653 : AOI221_X1 port map( B1 => n18936, B2 => n11349, C1 => n18930, C2 => 
                           n11350, A => n11351, ZN => n11334);
   U6654 : AOI211_X1 port map( C1 => registers_4_4_port, C2 => n18978, A => 
                           n11345, B => n11346, ZN => n11335);
   U6655 : NAND4_X1 port map( A1 => n11265, A2 => n11266, A3 => n11267, A4 => 
                           n11268, ZN => n7043);
   U6656 : AOI222_X1 port map( A1 => out_to_mem_5_port, A2 => n18917, B1 => 
                           n18909, B2 => n18203, C1 => registers_3_5_port, C2 
                           => n18903, ZN => n11265);
   U6657 : AOI221_X1 port map( B1 => n18936, B2 => n11282, C1 => n18930, C2 => 
                           n11283, A => n11284, ZN => n11266);
   U6658 : AOI211_X1 port map( C1 => registers_4_5_port, C2 => n18978, A => 
                           n11277, B => n11279, ZN => n11267);
   U6659 : NAND4_X1 port map( A1 => n11198, A2 => n11199, A3 => n11200, A4 => 
                           n11201, ZN => n7047);
   U6660 : AOI222_X1 port map( A1 => out_to_mem_6_port, A2 => n18917, B1 => 
                           n18909, B2 => n18204, C1 => registers_3_6_port, C2 
                           => n18903, ZN => n11198);
   U6661 : AOI221_X1 port map( B1 => n18936, B2 => n11214, C1 => n18930, C2 => 
                           n11215, A => n11216, ZN => n11199);
   U6662 : AOI211_X1 port map( C1 => registers_4_6_port, C2 => n18978, A => 
                           n11210, B => n11211, ZN => n11200);
   U6663 : NAND4_X1 port map( A1 => n11131, A2 => n11132, A3 => n11133, A4 => 
                           n11134, ZN => n7051);
   U6664 : AOI222_X1 port map( A1 => out_to_mem_7_port, A2 => n18917, B1 => 
                           n18909, B2 => n18205, C1 => registers_3_7_port, C2 
                           => n18903, ZN => n11131);
   U6665 : AOI221_X1 port map( B1 => n18936, B2 => n11147, C1 => n18930, C2 => 
                           n11148, A => n11149, ZN => n11132);
   U6666 : AOI211_X1 port map( C1 => registers_4_7_port, C2 => n18978, A => 
                           n11143, B => n11144, ZN => n11133);
   U6667 : NAND4_X1 port map( A1 => n11063, A2 => n11064, A3 => n11065, A4 => 
                           n11067, ZN => n7055);
   U6668 : AOI222_X1 port map( A1 => out_to_mem_8_port, A2 => n18917, B1 => 
                           n18909, B2 => n18206, C1 => registers_3_8_port, C2 
                           => n18903, ZN => n11063);
   U6669 : AOI221_X1 port map( B1 => n18936, B2 => n11080, C1 => n18930, C2 => 
                           n11081, A => n11082, ZN => n11064);
   U6670 : AOI211_X1 port map( C1 => registers_4_8_port, C2 => n18978, A => 
                           n11076, B => n11077, ZN => n11065);
   U6671 : NAND4_X1 port map( A1 => n10996, A2 => n10997, A3 => n10998, A4 => 
                           n10999, ZN => n7059);
   U6672 : AOI222_X1 port map( A1 => out_to_mem_9_port, A2 => n18917, B1 => 
                           n18909, B2 => n18207, C1 => registers_3_9_port, C2 
                           => n18903, ZN => n10996);
   U6673 : AOI221_X1 port map( B1 => n18936, B2 => n11012, C1 => n18930, C2 => 
                           n11014, A => n11015, ZN => n10997);
   U6674 : AOI211_X1 port map( C1 => registers_4_9_port, C2 => n18978, A => 
                           n11008, B => n11009, ZN => n10998);
   U6675 : NAND4_X1 port map( A1 => n10929, A2 => n10930, A3 => n10931, A4 => 
                           n10932, ZN => n7063);
   U6676 : AOI222_X1 port map( A1 => out_to_mem_10_port, A2 => n18917, B1 => 
                           n18909, B2 => n18208, C1 => registers_3_10_port, C2 
                           => n18903, ZN => n10929);
   U6677 : AOI221_X1 port map( B1 => n18936, B2 => n10945, C1 => n18930, C2 => 
                           n10946, A => n10947, ZN => n10930);
   U6678 : AOI211_X1 port map( C1 => registers_4_10_port, C2 => n18978, A => 
                           n10941, B => n10942, ZN => n10931);
   U6679 : NAND4_X1 port map( A1 => n10862, A2 => n10863, A3 => n10864, A4 => 
                           n10865, ZN => n7067);
   U6680 : AOI222_X1 port map( A1 => out_to_mem_11_port, A2 => n18917, B1 => 
                           n18909, B2 => n18209, C1 => registers_3_11_port, C2 
                           => n18903, ZN => n10862);
   U6681 : AOI221_X1 port map( B1 => n18936, B2 => n10878, C1 => n18930, C2 => 
                           n10879, A => n10880, ZN => n10863);
   U6682 : AOI211_X1 port map( C1 => registers_4_11_port, C2 => n18978, A => 
                           n10874, B => n10875, ZN => n10864);
   U6683 : NAND4_X1 port map( A1 => n10794, A2 => n10795, A3 => n10796, A4 => 
                           n10797, ZN => n7071);
   U6684 : AOI222_X1 port map( A1 => out_to_mem_12_port, A2 => n18917, B1 => 
                           n18910, B2 => n18210, C1 => registers_3_12_port, C2 
                           => n18904, ZN => n10794);
   U6685 : AOI221_X1 port map( B1 => n18937, B2 => n10811, C1 => n18931, C2 => 
                           n10812, A => n10813, ZN => n10795);
   U6686 : AOI211_X1 port map( C1 => registers_4_12_port, C2 => n18979, A => 
                           n10807, B => n10808, ZN => n10796);
   U6687 : NAND4_X1 port map( A1 => n10727, A2 => n10728, A3 => n10729, A4 => 
                           n10730, ZN => n7075);
   U6688 : AOI222_X1 port map( A1 => out_to_mem_13_port, A2 => n18917, B1 => 
                           n18910, B2 => n18211, C1 => registers_3_13_port, C2 
                           => n18904, ZN => n10727);
   U6689 : AOI221_X1 port map( B1 => n18937, B2 => n10743, C1 => n18931, C2 => 
                           n10744, A => n10745, ZN => n10728);
   U6690 : AOI211_X1 port map( C1 => registers_4_13_port, C2 => n18979, A => 
                           n10739, B => n10740, ZN => n10729);
   U6691 : NAND4_X1 port map( A1 => n10660, A2 => n10661, A3 => n10662, A4 => 
                           n10663, ZN => n7079);
   U6692 : AOI222_X1 port map( A1 => out_to_mem_14_port, A2 => n18917, B1 => 
                           n18910, B2 => n18212, C1 => registers_3_14_port, C2 
                           => n18904, ZN => n10660);
   U6693 : AOI221_X1 port map( B1 => n18937, B2 => n10676, C1 => n18931, C2 => 
                           n10677, A => n10678, ZN => n10661);
   U6694 : AOI211_X1 port map( C1 => registers_4_14_port, C2 => n18979, A => 
                           n10672, B => n10673, ZN => n10662);
   U6695 : NAND4_X1 port map( A1 => n10593, A2 => n10594, A3 => n10595, A4 => 
                           n10596, ZN => n7083);
   U6696 : AOI222_X1 port map( A1 => out_to_mem_15_port, A2 => n18917, B1 => 
                           n18910, B2 => n18213, C1 => registers_3_15_port, C2 
                           => n18904, ZN => n10593);
   U6697 : AOI221_X1 port map( B1 => n18937, B2 => n10609, C1 => n18931, C2 => 
                           n10610, A => n10611, ZN => n10594);
   U6698 : AOI211_X1 port map( C1 => registers_4_15_port, C2 => n18979, A => 
                           n10605, B => n10606, ZN => n10595);
   U6699 : NAND4_X1 port map( A1 => n10525, A2 => n10526, A3 => n10527, A4 => 
                           n10528, ZN => n7087);
   U6700 : AOI222_X1 port map( A1 => out_to_mem_16_port, A2 => n18917, B1 => 
                           n18910, B2 => n18214, C1 => registers_3_16_port, C2 
                           => n18904, ZN => n10525);
   U6701 : AOI221_X1 port map( B1 => n18937, B2 => n10542, C1 => n18931, C2 => 
                           n10543, A => n10544, ZN => n10526);
   U6702 : AOI211_X1 port map( C1 => registers_4_16_port, C2 => n18979, A => 
                           n10538, B => n10539, ZN => n10527);
   U6703 : NAND4_X1 port map( A1 => n10458, A2 => n10459, A3 => n10460, A4 => 
                           n10461, ZN => n7091);
   U6704 : AOI222_X1 port map( A1 => out_to_mem_17_port, A2 => n18917, B1 => 
                           n18910, B2 => n18215, C1 => registers_3_17_port, C2 
                           => n18904, ZN => n10458);
   U6705 : AOI221_X1 port map( B1 => n18937, B2 => n10474, C1 => n18931, C2 => 
                           n10475, A => n10476, ZN => n10459);
   U6706 : AOI211_X1 port map( C1 => registers_4_17_port, C2 => n18979, A => 
                           n10470, B => n10471, ZN => n10460);
   U6707 : NAND4_X1 port map( A1 => n10391, A2 => n10392, A3 => n10393, A4 => 
                           n10394, ZN => n7095);
   U6708 : AOI222_X1 port map( A1 => out_to_mem_18_port, A2 => n18917, B1 => 
                           n18910, B2 => n18216, C1 => registers_3_18_port, C2 
                           => n18904, ZN => n10391);
   U6709 : AOI221_X1 port map( B1 => n18937, B2 => n10407, C1 => n18931, C2 => 
                           n10408, A => n10409, ZN => n10392);
   U6710 : AOI211_X1 port map( C1 => registers_4_18_port, C2 => n18979, A => 
                           n10403, B => n10404, ZN => n10393);
   U6711 : NAND4_X1 port map( A1 => n10323, A2 => n10325, A3 => n10326, A4 => 
                           n10327, ZN => n7099);
   U6712 : AOI222_X1 port map( A1 => out_to_mem_19_port, A2 => n18916, B1 => 
                           n18910, B2 => n18217, C1 => registers_3_19_port, C2 
                           => n18904, ZN => n10323);
   U6713 : AOI221_X1 port map( B1 => n18937, B2 => n10340, C1 => n18931, C2 => 
                           n10341, A => n10342, ZN => n10325);
   U6714 : AOI211_X1 port map( C1 => registers_4_19_port, C2 => n18979, A => 
                           n10336, B => n10337, ZN => n10326);
   U6715 : NAND4_X1 port map( A1 => n10256, A2 => n10257, A3 => n10258, A4 => 
                           n10259, ZN => n7103);
   U6716 : AOI222_X1 port map( A1 => out_to_mem_20_port, A2 => n18916, B1 => 
                           n18910, B2 => n18218, C1 => registers_3_20_port, C2 
                           => n18904, ZN => n10256);
   U6717 : AOI221_X1 port map( B1 => n18937, B2 => n10273, C1 => n18931, C2 => 
                           n10274, A => n10275, ZN => n10257);
   U6718 : AOI211_X1 port map( C1 => registers_4_20_port, C2 => n18979, A => 
                           n10268, B => n10269, ZN => n10258);
   U6719 : NAND4_X1 port map( A1 => n10189, A2 => n10190, A3 => n10191, A4 => 
                           n10192, ZN => n7107);
   U6720 : AOI222_X1 port map( A1 => out_to_mem_21_port, A2 => n18916, B1 => 
                           n18910, B2 => n18219, C1 => registers_3_21_port, C2 
                           => n18904, ZN => n10189);
   U6721 : AOI221_X1 port map( B1 => n18937, B2 => n10205, C1 => n18931, C2 => 
                           n10206, A => n10207, ZN => n10190);
   U6722 : AOI211_X1 port map( C1 => registers_4_21_port, C2 => n18979, A => 
                           n10201, B => n10202, ZN => n10191);
   U6723 : NAND4_X1 port map( A1 => n10122, A2 => n10123, A3 => n10124, A4 => 
                           n10125, ZN => n7111);
   U6724 : AOI222_X1 port map( A1 => out_to_mem_22_port, A2 => n18916, B1 => 
                           n18910, B2 => n18220, C1 => registers_3_22_port, C2 
                           => n18904, ZN => n10122);
   U6725 : AOI221_X1 port map( B1 => n18937, B2 => n10138, C1 => n18931, C2 => 
                           n10139, A => n10140, ZN => n10123);
   U6726 : AOI211_X1 port map( C1 => registers_4_22_port, C2 => n18979, A => 
                           n10134, B => n10135, ZN => n10124);
   U6727 : NAND4_X1 port map( A1 => n10054, A2 => n10055, A3 => n10056, A4 => 
                           n10057, ZN => n7115);
   U6728 : AOI222_X1 port map( A1 => out_to_mem_23_port, A2 => n18916, B1 => 
                           n18910, B2 => n18221, C1 => registers_3_23_port, C2 
                           => n18904, ZN => n10054);
   U6729 : AOI221_X1 port map( B1 => n18937, B2 => n10071, C1 => n18931, C2 => 
                           n10072, A => n10073, ZN => n10055);
   U6730 : AOI211_X1 port map( C1 => registers_4_23_port, C2 => n18979, A => 
                           n10067, B => n10068, ZN => n10056);
   U6731 : NAND4_X1 port map( A1 => n9987, A2 => n9988, A3 => n9989, A4 => 
                           n9990, ZN => n7119);
   U6732 : AOI222_X1 port map( A1 => out_to_mem_24_port, A2 => n18916, B1 => 
                           n18911, B2 => n18222, C1 => registers_3_24_port, C2 
                           => n18905, ZN => n9987);
   U6733 : AOI221_X1 port map( B1 => n18938, B2 => n10003, C1 => n18932, C2 => 
                           n10004, A => n10005, ZN => n9988);
   U6734 : AOI211_X1 port map( C1 => registers_4_24_port, C2 => n18980, A => 
                           n9999, B => n10000, ZN => n9989);
   U6735 : NAND4_X1 port map( A1 => n9920, A2 => n9921, A3 => n9922, A4 => 
                           n9923, ZN => n7123);
   U6736 : AOI222_X1 port map( A1 => out_to_mem_25_port, A2 => n18916, B1 => 
                           n18911, B2 => n18223, C1 => registers_3_25_port, C2 
                           => n18905, ZN => n9920);
   U6737 : AOI221_X1 port map( B1 => n18938, B2 => n9936, C1 => n18932, C2 => 
                           n9937, A => n9938, ZN => n9921);
   U6738 : AOI211_X1 port map( C1 => registers_4_25_port, C2 => n18980, A => 
                           n9932, B => n9933, ZN => n9922);
   U6739 : NAND4_X1 port map( A1 => n9853, A2 => n9854, A3 => n9855, A4 => 
                           n9856, ZN => n7127);
   U6740 : AOI222_X1 port map( A1 => out_to_mem_26_port, A2 => n18916, B1 => 
                           n18911, B2 => n18224, C1 => registers_3_26_port, C2 
                           => n18905, ZN => n9853);
   U6741 : AOI221_X1 port map( B1 => n18938, B2 => n9869, C1 => n18932, C2 => 
                           n9870, A => n9871, ZN => n9854);
   U6742 : AOI211_X1 port map( C1 => registers_4_26_port, C2 => n18980, A => 
                           n9865, B => n9866, ZN => n9855);
   U6743 : NAND4_X1 port map( A1 => n9785, A2 => n9786, A3 => n9787, A4 => 
                           n9788, ZN => n7131);
   U6744 : AOI222_X1 port map( A1 => out_to_mem_27_port, A2 => n18916, B1 => 
                           n18911, B2 => n18225, C1 => registers_3_27_port, C2 
                           => n18905, ZN => n9785);
   U6745 : AOI221_X1 port map( B1 => n18938, B2 => n9802, C1 => n18932, C2 => 
                           n9803, A => n9804, ZN => n9786);
   U6746 : AOI211_X1 port map( C1 => registers_4_27_port, C2 => n18980, A => 
                           n9798, B => n9799, ZN => n9787);
   U6747 : NAND4_X1 port map( A1 => n9718, A2 => n9719, A3 => n9720, A4 => 
                           n9721, ZN => n7135);
   U6748 : AOI222_X1 port map( A1 => out_to_mem_28_port, A2 => n18916, B1 => 
                           n18911, B2 => n18226, C1 => registers_3_28_port, C2 
                           => n18905, ZN => n9718);
   U6749 : AOI221_X1 port map( B1 => n18938, B2 => n9734, C1 => n18932, C2 => 
                           n9735, A => n9736, ZN => n9719);
   U6750 : AOI211_X1 port map( C1 => registers_4_28_port, C2 => n18980, A => 
                           n9730, B => n9731, ZN => n9720);
   U6751 : NAND4_X1 port map( A1 => n9651, A2 => n9652, A3 => n9653, A4 => 
                           n9654, ZN => n7139);
   U6752 : AOI222_X1 port map( A1 => out_to_mem_29_port, A2 => n18916, B1 => 
                           n18911, B2 => n18227, C1 => registers_3_29_port, C2 
                           => n18905, ZN => n9651);
   U6753 : AOI221_X1 port map( B1 => n18938, B2 => n9667, C1 => n18932, C2 => 
                           n9668, A => n9669, ZN => n9652);
   U6754 : AOI211_X1 port map( C1 => registers_4_29_port, C2 => n18980, A => 
                           n9663, B => n9664, ZN => n9653);
   U6755 : NAND4_X1 port map( A1 => n9584, A2 => n9585, A3 => n9586, A4 => 
                           n9587, ZN => n7143);
   U6756 : AOI222_X1 port map( A1 => out_to_mem_30_port, A2 => n18916, B1 => 
                           n18911, B2 => n18228, C1 => registers_3_30_port, C2 
                           => n18905, ZN => n9584);
   U6757 : AOI221_X1 port map( B1 => n18938, B2 => n9600, C1 => n18932, C2 => 
                           n9601, A => n9602, ZN => n9585);
   U6758 : AOI211_X1 port map( C1 => registers_4_30_port, C2 => n18980, A => 
                           n9596, B => n9597, ZN => n9586);
   U6759 : NAND4_X1 port map( A1 => n9516, A2 => n9517, A3 => n9518, A4 => 
                           n9519, ZN => n7147);
   U6760 : AOI222_X1 port map( A1 => out_to_mem_31_port, A2 => n18916, B1 => 
                           n18911, B2 => n18229, C1 => registers_3_31_port, C2 
                           => n18905, ZN => n9516);
   U6761 : AOI221_X1 port map( B1 => n18938, B2 => n9533, C1 => n18932, C2 => 
                           n9534, A => n9535, ZN => n9517);
   U6762 : AOI211_X1 port map( C1 => registers_4_31_port, C2 => n18980, A => 
                           n9528, B => n9529, ZN => n9518);
   U6763 : NAND4_X1 port map( A1 => n9449, A2 => n9450, A3 => n9451, A4 => 
                           n9452, ZN => n7151);
   U6764 : AOI222_X1 port map( A1 => out_to_mem_32_port, A2 => n18916, B1 => 
                           n18911, B2 => n18230, C1 => registers_3_32_port, C2 
                           => n18905, ZN => n9449);
   U6765 : AOI221_X1 port map( B1 => n18938, B2 => n9465, C1 => n18932, C2 => 
                           n9466, A => n9467, ZN => n9450);
   U6766 : AOI211_X1 port map( C1 => registers_4_32_port, C2 => n18980, A => 
                           n9461, B => n9462, ZN => n9451);
   U6767 : NAND4_X1 port map( A1 => n9382, A2 => n9383, A3 => n9384, A4 => 
                           n9385, ZN => n7155);
   U6768 : AOI222_X1 port map( A1 => out_to_mem_33_port, A2 => n18915, B1 => 
                           n18911, B2 => n18231, C1 => registers_3_33_port, C2 
                           => n18905, ZN => n9382);
   U6769 : AOI221_X1 port map( B1 => n18938, B2 => n9398, C1 => n18932, C2 => 
                           n9399, A => n9400, ZN => n9383);
   U6770 : AOI211_X1 port map( C1 => registers_4_33_port, C2 => n18980, A => 
                           n9394, B => n9395, ZN => n9384);
   U6771 : NAND4_X1 port map( A1 => n9314, A2 => n9315, A3 => n9316, A4 => 
                           n9317, ZN => n7159);
   U6772 : AOI222_X1 port map( A1 => out_to_mem_34_port, A2 => n18915, B1 => 
                           n18911, B2 => n18232, C1 => registers_3_34_port, C2 
                           => n18905, ZN => n9314);
   U6773 : AOI221_X1 port map( B1 => n18938, B2 => n9331, C1 => n18932, C2 => 
                           n9332, A => n9333, ZN => n9315);
   U6774 : AOI211_X1 port map( C1 => registers_4_34_port, C2 => n18980, A => 
                           n9327, B => n9328, ZN => n9316);
   U6775 : NAND4_X1 port map( A1 => n7007, A2 => n7008, A3 => n7009, A4 => 
                           n7010, ZN => n7163);
   U6776 : AOI222_X1 port map( A1 => out_to_mem_35_port, A2 => n18915, B1 => 
                           n18911, B2 => n18233, C1 => registers_3_35_port, C2 
                           => n18905, ZN => n7007);
   U6777 : AOI221_X1 port map( B1 => n18938, B2 => n9263, C1 => n18932, C2 => 
                           n9264, A => n9266, ZN => n7008);
   U6778 : AOI211_X1 port map( C1 => registers_4_35_port, C2 => n18980, A => 
                           n7019, B => n7020, ZN => n7009);
   U6779 : NAND4_X1 port map( A1 => n6940, A2 => n6941, A3 => n6942, A4 => 
                           n6943, ZN => n7167);
   U6780 : AOI222_X1 port map( A1 => out_to_mem_36_port, A2 => n18916, B1 => 
                           n18912, B2 => n18234, C1 => registers_3_36_port, C2 
                           => n18906, ZN => n6940);
   U6781 : AOI221_X1 port map( B1 => n18939, B2 => n6957, C1 => n18933, C2 => 
                           n6958, A => n6959, ZN => n6941);
   U6782 : AOI211_X1 port map( C1 => registers_4_36_port, C2 => n18981, A => 
                           n6953, B => n6954, ZN => n6942);
   U6783 : NAND4_X1 port map( A1 => n6874, A2 => n6875, A3 => n6876, A4 => 
                           n6877, ZN => n7171);
   U6784 : AOI222_X1 port map( A1 => out_to_mem_37_port, A2 => n18917, B1 => 
                           n18912, B2 => n18235, C1 => registers_3_37_port, C2 
                           => n18906, ZN => n6874);
   U6785 : AOI221_X1 port map( B1 => n18939, B2 => n6890, C1 => n18933, C2 => 
                           n6891, A => n6892, ZN => n6875);
   U6786 : AOI211_X1 port map( C1 => registers_4_37_port, C2 => n18981, A => 
                           n6886, B => n6887, ZN => n6876);
   U6787 : AND3_X1 port map( A1 => count3(0), A2 => n11672, A3 => n11688, ZN =>
                           n11673);
   U6788 : AOI21_X1 port map( B1 => count3(2), B2 => count3(1), A => n11747, ZN
                           => n11746);
   U6789 : NAND4_X1 port map( A1 => n11624, A2 => n11625, A3 => n11626, A4 => 
                           n11627, ZN => n7024);
   U6790 : AOI221_X1 port map( B1 => n19092, B2 => n11618, C1 => n19086, C2 => 
                           n11619, A => n11659, ZN => n11624);
   U6791 : AOI221_X1 port map( B1 => n19116, B2 => registers_15_0_port, C1 => 
                           n19110, C2 => registers_14_0_port, A => n11657, ZN 
                           => n11625);
   U6792 : NOR4_X1 port map( A1 => n11647, A2 => n11649, A3 => n11650, A4 => 
                           n11651, ZN => n11626);
   U6793 : NAND4_X1 port map( A1 => n11576, A2 => n11577, A3 => n11578, A4 => 
                           n11579, ZN => n7025);
   U6794 : AOI221_X1 port map( B1 => n19291, B2 => n11618, C1 => n19285, C2 => 
                           n11619, A => n11620, ZN => n11576);
   U6795 : NOR4_X1 port map( A1 => n11607, A2 => n11608, A3 => n11609, A4 => 
                           n11610, ZN => n11578);
   U6796 : AOI221_X1 port map( B1 => n19315, B2 => registers_15_0_port, C1 => 
                           n19309, C2 => registers_14_0_port, A => n11615, ZN 
                           => n11577);
   U6797 : NAND4_X1 port map( A1 => n11516, A2 => n11517, A3 => n11518, A4 => 
                           n11519, ZN => n7028);
   U6798 : AOI221_X1 port map( B1 => n19092, B2 => n11513, C1 => n19086, C2 => 
                           n11514, A => n11533, ZN => n11516);
   U6799 : AOI221_X1 port map( B1 => n19116, B2 => registers_15_1_port, C1 => 
                           n19110, C2 => registers_14_1_port, A => n11532, ZN 
                           => n11517);
   U6800 : NOR4_X1 port map( A1 => n11528, A2 => n11529, A3 => n11530, A4 => 
                           n11531, ZN => n11518);
   U6801 : NAND4_X1 port map( A1 => n11488, A2 => n11490, A3 => n11491, A4 => 
                           n11492, ZN => n7029);
   U6802 : AOI221_X1 port map( B1 => n19291, B2 => n11513, C1 => n19285, C2 => 
                           n11514, A => n11515, ZN => n11488);
   U6803 : NOR4_X1 port map( A1 => n11508, A2 => n11509, A3 => n11510, A4 => 
                           n11511, ZN => n11491);
   U6804 : AOI221_X1 port map( B1 => n19315, B2 => registers_15_1_port, C1 => 
                           n19309, C2 => registers_14_1_port, A => n11512, ZN 
                           => n11490);
   U6805 : NAND4_X1 port map( A1 => n11449, A2 => n11450, A3 => n11451, A4 => 
                           n11452, ZN => n7032);
   U6806 : AOI221_X1 port map( B1 => n19092, B2 => n11446, C1 => n19086, C2 => 
                           n11447, A => n11466, ZN => n11449);
   U6807 : AOI221_X1 port map( B1 => n19116, B2 => registers_15_2_port, C1 => 
                           n19110, C2 => registers_14_2_port, A => n11465, ZN 
                           => n11450);
   U6808 : NOR4_X1 port map( A1 => n11461, A2 => n11462, A3 => n11463, A4 => 
                           n11464, ZN => n11451);
   U6809 : NAND4_X1 port map( A1 => n11421, A2 => n11422, A3 => n11423, A4 => 
                           n11424, ZN => n7033);
   U6810 : AOI221_X1 port map( B1 => n19291, B2 => n11446, C1 => n19285, C2 => 
                           n11447, A => n11448, ZN => n11421);
   U6811 : NOR4_X1 port map( A1 => n11441, A2 => n11442, A3 => n11443, A4 => 
                           n11444, ZN => n11423);
   U6812 : AOI221_X1 port map( B1 => n19315, B2 => registers_15_2_port, C1 => 
                           n19309, C2 => registers_14_2_port, A => n11445, ZN 
                           => n11422);
   U6813 : NAND4_X1 port map( A1 => n11381, A2 => n11382, A3 => n11383, A4 => 
                           n11385, ZN => n7036);
   U6814 : AOI221_X1 port map( B1 => n19092, B2 => n11378, C1 => n19086, C2 => 
                           n11379, A => n11399, ZN => n11381);
   U6815 : AOI221_X1 port map( B1 => n19116, B2 => registers_15_3_port, C1 => 
                           n19110, C2 => registers_14_3_port, A => n11398, ZN 
                           => n11382);
   U6816 : NOR4_X1 port map( A1 => n11394, A2 => n11395, A3 => n11396, A4 => 
                           n11397, ZN => n11383);
   U6817 : NAND4_X1 port map( A1 => n11354, A2 => n11355, A3 => n11356, A4 => 
                           n11357, ZN => n7037);
   U6818 : AOI221_X1 port map( B1 => n19291, B2 => n11378, C1 => n19285, C2 => 
                           n11379, A => n11380, ZN => n11354);
   U6819 : NOR4_X1 port map( A1 => n11373, A2 => n11374, A3 => n11375, A4 => 
                           n11376, ZN => n11356);
   U6820 : AOI221_X1 port map( B1 => n19315, B2 => registers_15_3_port, C1 => 
                           n19309, C2 => registers_14_3_port, A => n11377, ZN 
                           => n11355);
   U6821 : NAND4_X1 port map( A1 => n11314, A2 => n11315, A3 => n11316, A4 => 
                           n11317, ZN => n7040);
   U6822 : AOI221_X1 port map( B1 => n19092, B2 => n11311, C1 => n19086, C2 => 
                           n11312, A => n11332, ZN => n11314);
   U6823 : AOI221_X1 port map( B1 => n19116, B2 => registers_15_4_port, C1 => 
                           n19110, C2 => registers_14_4_port, A => n11330, ZN 
                           => n11315);
   U6824 : NOR4_X1 port map( A1 => n11326, A2 => n11327, A3 => n11328, A4 => 
                           n11329, ZN => n11316);
   U6825 : NAND4_X1 port map( A1 => n11287, A2 => n11288, A3 => n11289, A4 => 
                           n11290, ZN => n7041);
   U6826 : AOI221_X1 port map( B1 => n19291, B2 => n11311, C1 => n19285, C2 => 
                           n11312, A => n11313, ZN => n11287);
   U6827 : NOR4_X1 port map( A1 => n11306, A2 => n11307, A3 => n11308, A4 => 
                           n11309, ZN => n11289);
   U6828 : AOI221_X1 port map( B1 => n19315, B2 => registers_15_4_port, C1 => 
                           n19309, C2 => registers_14_4_port, A => n11310, ZN 
                           => n11288);
   U6829 : NAND4_X1 port map( A1 => n11247, A2 => n11248, A3 => n11249, A4 => 
                           n11250, ZN => n7044);
   U6830 : AOI221_X1 port map( B1 => n19092, B2 => n11244, C1 => n19086, C2 => 
                           n11245, A => n11264, ZN => n11247);
   U6831 : AOI221_X1 port map( B1 => n19116, B2 => registers_15_5_port, C1 => 
                           n19110, C2 => registers_14_5_port, A => n11263, ZN 
                           => n11248);
   U6832 : NOR4_X1 port map( A1 => n11259, A2 => n11260, A3 => n11261, A4 => 
                           n11262, ZN => n11249);
   U6833 : NAND4_X1 port map( A1 => n11219, A2 => n11220, A3 => n11221, A4 => 
                           n11222, ZN => n7045);
   U6834 : AOI221_X1 port map( B1 => n19291, B2 => n11244, C1 => n19285, C2 => 
                           n11245, A => n11246, ZN => n11219);
   U6835 : NOR4_X1 port map( A1 => n11239, A2 => n11240, A3 => n11241, A4 => 
                           n11242, ZN => n11221);
   U6836 : AOI221_X1 port map( B1 => n19315, B2 => registers_15_5_port, C1 => 
                           n19309, C2 => registers_14_5_port, A => n11243, ZN 
                           => n11220);
   U6837 : NAND4_X1 port map( A1 => n11180, A2 => n11181, A3 => n11182, A4 => 
                           n11183, ZN => n7048);
   U6838 : AOI221_X1 port map( B1 => n19092, B2 => n11177, C1 => n19086, C2 => 
                           n11178, A => n11197, ZN => n11180);
   U6839 : AOI221_X1 port map( B1 => n19116, B2 => registers_15_6_port, C1 => 
                           n19110, C2 => registers_14_6_port, A => n11196, ZN 
                           => n11181);
   U6840 : NOR4_X1 port map( A1 => n11192, A2 => n11193, A3 => n11194, A4 => 
                           n11195, ZN => n11182);
   U6841 : NAND4_X1 port map( A1 => n11152, A2 => n11153, A3 => n11154, A4 => 
                           n11155, ZN => n7049);
   U6842 : AOI221_X1 port map( B1 => n19291, B2 => n11177, C1 => n19285, C2 => 
                           n11178, A => n11179, ZN => n11152);
   U6843 : NOR4_X1 port map( A1 => n11171, A2 => n11173, A3 => n11174, A4 => 
                           n11175, ZN => n11154);
   U6844 : AOI221_X1 port map( B1 => n19315, B2 => registers_15_6_port, C1 => 
                           n19309, C2 => registers_14_6_port, A => n11176, ZN 
                           => n11153);
   U6845 : NAND4_X1 port map( A1 => n11112, A2 => n11113, A3 => n11114, A4 => 
                           n11115, ZN => n7052);
   U6846 : AOI221_X1 port map( B1 => n19092, B2 => n11109, C1 => n19086, C2 => 
                           n11110, A => n11130, ZN => n11112);
   U6847 : AOI221_X1 port map( B1 => n19116, B2 => registers_15_7_port, C1 => 
                           n19110, C2 => registers_14_7_port, A => n11129, ZN 
                           => n11113);
   U6848 : NOR4_X1 port map( A1 => n11125, A2 => n11126, A3 => n11127, A4 => 
                           n11128, ZN => n11114);
   U6849 : NAND4_X1 port map( A1 => n11085, A2 => n11086, A3 => n11087, A4 => 
                           n11088, ZN => n7053);
   U6850 : AOI221_X1 port map( B1 => n19291, B2 => n11109, C1 => n19285, C2 => 
                           n11110, A => n11111, ZN => n11085);
   U6851 : NOR4_X1 port map( A1 => n11104, A2 => n11105, A3 => n11106, A4 => 
                           n11107, ZN => n11087);
   U6852 : AOI221_X1 port map( B1 => n19315, B2 => registers_15_7_port, C1 => 
                           n19309, C2 => registers_14_7_port, A => n11108, ZN 
                           => n11086);
   U6853 : NAND4_X1 port map( A1 => n11045, A2 => n11046, A3 => n11047, A4 => 
                           n11048, ZN => n7056);
   U6854 : AOI221_X1 port map( B1 => n19092, B2 => n11042, C1 => n19086, C2 => 
                           n11043, A => n11062, ZN => n11045);
   U6855 : AOI221_X1 port map( B1 => n19116, B2 => registers_15_8_port, C1 => 
                           n19110, C2 => registers_14_8_port, A => n11061, ZN 
                           => n11046);
   U6856 : NOR4_X1 port map( A1 => n11057, A2 => n11058, A3 => n11059, A4 => 
                           n11060, ZN => n11047);
   U6857 : NAND4_X1 port map( A1 => n11018, A2 => n11019, A3 => n11020, A4 => 
                           n11021, ZN => n7057);
   U6858 : AOI221_X1 port map( B1 => n19291, B2 => n11042, C1 => n19285, C2 => 
                           n11043, A => n11044, ZN => n11018);
   U6859 : NOR4_X1 port map( A1 => n11037, A2 => n11038, A3 => n11039, A4 => 
                           n11040, ZN => n11020);
   U6860 : AOI221_X1 port map( B1 => n19315, B2 => registers_15_8_port, C1 => 
                           n19309, C2 => registers_14_8_port, A => n11041, ZN 
                           => n11019);
   U6861 : NAND4_X1 port map( A1 => n10978, A2 => n10979, A3 => n10980, A4 => 
                           n10981, ZN => n7060);
   U6862 : AOI221_X1 port map( B1 => n19092, B2 => n10975, C1 => n19086, C2 => 
                           n10976, A => n10995, ZN => n10978);
   U6863 : AOI221_X1 port map( B1 => n19116, B2 => registers_15_9_port, C1 => 
                           n19110, C2 => registers_14_9_port, A => n10994, ZN 
                           => n10979);
   U6864 : NOR4_X1 port map( A1 => n10990, A2 => n10991, A3 => n10992, A4 => 
                           n10993, ZN => n10980);
   U6865 : NAND4_X1 port map( A1 => n10950, A2 => n10951, A3 => n10952, A4 => 
                           n10953, ZN => n7061);
   U6866 : AOI221_X1 port map( B1 => n19291, B2 => n10975, C1 => n19285, C2 => 
                           n10976, A => n10977, ZN => n10950);
   U6867 : NOR4_X1 port map( A1 => n10970, A2 => n10971, A3 => n10972, A4 => 
                           n10973, ZN => n10952);
   U6868 : AOI221_X1 port map( B1 => n19315, B2 => registers_15_9_port, C1 => 
                           n19309, C2 => registers_14_9_port, A => n10974, ZN 
                           => n10951);
   U6869 : NAND4_X1 port map( A1 => n10911, A2 => n10912, A3 => n10913, A4 => 
                           n10914, ZN => n7064);
   U6870 : AOI221_X1 port map( B1 => n19092, B2 => n10908, C1 => n19086, C2 => 
                           n10909, A => n10928, ZN => n10911);
   U6871 : AOI221_X1 port map( B1 => n19116, B2 => registers_15_10_port, C1 => 
                           n19110, C2 => registers_14_10_port, A => n10927, ZN 
                           => n10912);
   U6872 : NOR4_X1 port map( A1 => n10923, A2 => n10924, A3 => n10925, A4 => 
                           n10926, ZN => n10913);
   U6873 : NAND4_X1 port map( A1 => n10883, A2 => n10884, A3 => n10885, A4 => 
                           n10886, ZN => n7065);
   U6874 : AOI221_X1 port map( B1 => n19291, B2 => n10908, C1 => n19285, C2 => 
                           n10909, A => n10910, ZN => n10883);
   U6875 : NOR4_X1 port map( A1 => n10902, A2 => n10903, A3 => n10904, A4 => 
                           n10905, ZN => n10885);
   U6876 : AOI221_X1 port map( B1 => n19315, B2 => registers_15_10_port, C1 => 
                           n19309, C2 => registers_14_10_port, A => n10906, ZN 
                           => n10884);
   U6877 : NAND4_X1 port map( A1 => n10843, A2 => n10844, A3 => n10845, A4 => 
                           n10846, ZN => n7068);
   U6878 : AOI221_X1 port map( B1 => n19092, B2 => n10840, C1 => n19086, C2 => 
                           n10841, A => n10861, ZN => n10843);
   U6879 : AOI221_X1 port map( B1 => n19116, B2 => registers_15_11_port, C1 => 
                           n19110, C2 => registers_14_11_port, A => n10860, ZN 
                           => n10844);
   U6880 : NOR4_X1 port map( A1 => n10856, A2 => n10857, A3 => n10858, A4 => 
                           n10859, ZN => n10845);
   U6881 : NAND4_X1 port map( A1 => n10816, A2 => n10817, A3 => n10818, A4 => 
                           n10819, ZN => n7069);
   U6882 : AOI221_X1 port map( B1 => n19291, B2 => n10840, C1 => n19285, C2 => 
                           n10841, A => n10842, ZN => n10816);
   U6883 : NOR4_X1 port map( A1 => n10835, A2 => n10836, A3 => n10837, A4 => 
                           n10838, ZN => n10818);
   U6884 : AOI221_X1 port map( B1 => n19315, B2 => registers_15_11_port, C1 => 
                           n19309, C2 => registers_14_11_port, A => n10839, ZN 
                           => n10817);
   U6885 : NAND4_X1 port map( A1 => n10776, A2 => n10777, A3 => n10778, A4 => 
                           n10779, ZN => n7072);
   U6886 : AOI221_X1 port map( B1 => n19093, B2 => n10773, C1 => n19087, C2 => 
                           n10774, A => n10793, ZN => n10776);
   U6887 : AOI221_X1 port map( B1 => n19117, B2 => registers_15_12_port, C1 => 
                           n19111, C2 => registers_14_12_port, A => n10792, ZN 
                           => n10777);
   U6888 : NOR4_X1 port map( A1 => n10788, A2 => n10789, A3 => n10790, A4 => 
                           n10791, ZN => n10778);
   U6889 : NAND4_X1 port map( A1 => n10749, A2 => n10750, A3 => n10751, A4 => 
                           n10752, ZN => n7073);
   U6890 : AOI221_X1 port map( B1 => n19292, B2 => n10773, C1 => n19286, C2 => 
                           n10774, A => n10775, ZN => n10749);
   U6891 : NOR4_X1 port map( A1 => n10768, A2 => n10769, A3 => n10770, A4 => 
                           n10771, ZN => n10751);
   U6892 : AOI221_X1 port map( B1 => n19316, B2 => registers_15_12_port, C1 => 
                           n19310, C2 => registers_14_12_port, A => n10772, ZN 
                           => n10750);
   U6893 : NAND4_X1 port map( A1 => n10709, A2 => n10710, A3 => n10711, A4 => 
                           n10712, ZN => n7076);
   U6894 : AOI221_X1 port map( B1 => n19093, B2 => n10706, C1 => n19087, C2 => 
                           n10707, A => n10726, ZN => n10709);
   U6895 : AOI221_X1 port map( B1 => n19117, B2 => registers_15_13_port, C1 => 
                           n19111, C2 => registers_14_13_port, A => n10725, ZN 
                           => n10710);
   U6896 : NOR4_X1 port map( A1 => n10721, A2 => n10722, A3 => n10723, A4 => 
                           n10724, ZN => n10711);
   U6897 : NAND4_X1 port map( A1 => n10681, A2 => n10682, A3 => n10683, A4 => 
                           n10684, ZN => n7077);
   U6898 : AOI221_X1 port map( B1 => n19292, B2 => n10706, C1 => n19286, C2 => 
                           n10707, A => n10708, ZN => n10681);
   U6899 : NOR4_X1 port map( A1 => n10701, A2 => n10702, A3 => n10703, A4 => 
                           n10704, ZN => n10683);
   U6900 : AOI221_X1 port map( B1 => n19316, B2 => registers_15_13_port, C1 => 
                           n19310, C2 => registers_14_13_port, A => n10705, ZN 
                           => n10682);
   U6901 : NAND4_X1 port map( A1 => n10641, A2 => n10643, A3 => n10644, A4 => 
                           n10645, ZN => n7080);
   U6902 : AOI221_X1 port map( B1 => n19093, B2 => n10638, C1 => n19087, C2 => 
                           n10639, A => n10659, ZN => n10641);
   U6903 : AOI221_X1 port map( B1 => n19117, B2 => registers_15_14_port, C1 => 
                           n19111, C2 => registers_14_14_port, A => n10658, ZN 
                           => n10643);
   U6904 : NOR4_X1 port map( A1 => n10654, A2 => n10655, A3 => n10656, A4 => 
                           n10657, ZN => n10644);
   U6905 : NAND4_X1 port map( A1 => n10614, A2 => n10615, A3 => n10616, A4 => 
                           n10617, ZN => n7081);
   U6906 : AOI221_X1 port map( B1 => n19292, B2 => n10638, C1 => n19286, C2 => 
                           n10639, A => n10640, ZN => n10614);
   U6907 : NOR4_X1 port map( A1 => n10633, A2 => n10634, A3 => n10635, A4 => 
                           n10636, ZN => n10616);
   U6908 : AOI221_X1 port map( B1 => n19316, B2 => registers_15_14_port, C1 => 
                           n19310, C2 => registers_14_14_port, A => n10637, ZN 
                           => n10615);
   U6909 : NAND4_X1 port map( A1 => n10574, A2 => n10575, A3 => n10576, A4 => 
                           n10577, ZN => n7084);
   U6910 : AOI221_X1 port map( B1 => n19093, B2 => n10571, C1 => n19087, C2 => 
                           n10572, A => n10592, ZN => n10574);
   U6911 : AOI221_X1 port map( B1 => n19117, B2 => registers_15_15_port, C1 => 
                           n19111, C2 => registers_14_15_port, A => n10591, ZN 
                           => n10575);
   U6912 : NOR4_X1 port map( A1 => n10586, A2 => n10587, A3 => n10588, A4 => 
                           n10590, ZN => n10576);
   U6913 : NAND4_X1 port map( A1 => n10547, A2 => n10548, A3 => n10549, A4 => 
                           n10550, ZN => n7085);
   U6914 : AOI221_X1 port map( B1 => n19292, B2 => n10571, C1 => n19286, C2 => 
                           n10572, A => n10573, ZN => n10547);
   U6915 : NOR4_X1 port map( A1 => n10566, A2 => n10567, A3 => n10568, A4 => 
                           n10569, ZN => n10549);
   U6916 : AOI221_X1 port map( B1 => n19316, B2 => registers_15_15_port, C1 => 
                           n19310, C2 => registers_14_15_port, A => n10570, ZN 
                           => n10548);
   U6917 : NAND4_X1 port map( A1 => n10507, A2 => n10508, A3 => n10509, A4 => 
                           n10510, ZN => n7088);
   U6918 : AOI221_X1 port map( B1 => n19093, B2 => n10504, C1 => n19087, C2 => 
                           n10505, A => n10524, ZN => n10507);
   U6919 : AOI221_X1 port map( B1 => n19117, B2 => registers_15_16_port, C1 => 
                           n19111, C2 => registers_14_16_port, A => n10523, ZN 
                           => n10508);
   U6920 : NOR4_X1 port map( A1 => n10519, A2 => n10520, A3 => n10521, A4 => 
                           n10522, ZN => n10509);
   U6921 : NAND4_X1 port map( A1 => n10479, A2 => n10480, A3 => n10481, A4 => 
                           n10482, ZN => n7089);
   U6922 : AOI221_X1 port map( B1 => n19292, B2 => n10504, C1 => n19286, C2 => 
                           n10505, A => n10506, ZN => n10479);
   U6923 : NOR4_X1 port map( A1 => n10499, A2 => n10500, A3 => n10501, A4 => 
                           n10502, ZN => n10481);
   U6924 : AOI221_X1 port map( B1 => n19316, B2 => registers_15_16_port, C1 => 
                           n19310, C2 => registers_14_16_port, A => n10503, ZN 
                           => n10480);
   U6925 : NAND4_X1 port map( A1 => n10440, A2 => n10441, A3 => n10442, A4 => 
                           n10443, ZN => n7092);
   U6926 : AOI221_X1 port map( B1 => n19093, B2 => n10437, C1 => n19087, C2 => 
                           n10438, A => n10457, ZN => n10440);
   U6927 : AOI221_X1 port map( B1 => n19117, B2 => registers_15_17_port, C1 => 
                           n19111, C2 => registers_14_17_port, A => n10456, ZN 
                           => n10441);
   U6928 : NOR4_X1 port map( A1 => n10452, A2 => n10453, A3 => n10454, A4 => 
                           n10455, ZN => n10442);
   U6929 : NAND4_X1 port map( A1 => n10412, A2 => n10413, A3 => n10414, A4 => 
                           n10415, ZN => n7093);
   U6930 : AOI221_X1 port map( B1 => n19292, B2 => n10437, C1 => n19286, C2 => 
                           n10438, A => n10439, ZN => n10412);
   U6931 : NOR4_X1 port map( A1 => n10432, A2 => n10433, A3 => n10434, A4 => 
                           n10435, ZN => n10414);
   U6932 : AOI221_X1 port map( B1 => n19316, B2 => registers_15_17_port, C1 => 
                           n19310, C2 => registers_14_17_port, A => n10436, ZN 
                           => n10413);
   U6933 : NAND4_X1 port map( A1 => n10372, A2 => n10373, A3 => n10374, A4 => 
                           n10375, ZN => n7096);
   U6934 : AOI221_X1 port map( B1 => n19093, B2 => n10369, C1 => n19087, C2 => 
                           n10370, A => n10390, ZN => n10372);
   U6935 : AOI221_X1 port map( B1 => n19117, B2 => registers_15_18_port, C1 => 
                           n19111, C2 => registers_14_18_port, A => n10389, ZN 
                           => n10373);
   U6936 : NOR4_X1 port map( A1 => n10385, A2 => n10386, A3 => n10387, A4 => 
                           n10388, ZN => n10374);
   U6937 : NAND4_X1 port map( A1 => n10345, A2 => n10346, A3 => n10347, A4 => 
                           n10348, ZN => n7097);
   U6938 : AOI221_X1 port map( B1 => n19292, B2 => n10369, C1 => n19286, C2 => 
                           n10370, A => n10371, ZN => n10345);
   U6939 : NOR4_X1 port map( A1 => n10364, A2 => n10365, A3 => n10366, A4 => 
                           n10367, ZN => n10347);
   U6940 : AOI221_X1 port map( B1 => n19316, B2 => registers_15_18_port, C1 => 
                           n19310, C2 => registers_14_18_port, A => n10368, ZN 
                           => n10346);
   U6941 : NAND4_X1 port map( A1 => n10305, A2 => n10306, A3 => n10307, A4 => 
                           n10308, ZN => n7100);
   U6942 : AOI221_X1 port map( B1 => n19093, B2 => n10302, C1 => n19087, C2 => 
                           n10303, A => n10322, ZN => n10305);
   U6943 : AOI221_X1 port map( B1 => n19117, B2 => registers_15_19_port, C1 => 
                           n19111, C2 => registers_14_19_port, A => n10321, ZN 
                           => n10306);
   U6944 : NOR4_X1 port map( A1 => n10317, A2 => n10318, A3 => n10319, A4 => 
                           n10320, ZN => n10307);
   U6945 : NAND4_X1 port map( A1 => n10278, A2 => n10279, A3 => n10280, A4 => 
                           n10281, ZN => n7101);
   U6946 : AOI221_X1 port map( B1 => n19292, B2 => n10302, C1 => n19286, C2 => 
                           n10303, A => n10304, ZN => n10278);
   U6947 : NOR4_X1 port map( A1 => n10297, A2 => n10298, A3 => n10299, A4 => 
                           n10300, ZN => n10280);
   U6948 : AOI221_X1 port map( B1 => n19316, B2 => registers_15_19_port, C1 => 
                           n19310, C2 => registers_14_19_port, A => n10301, ZN 
                           => n10279);
   U6949 : NAND4_X1 port map( A1 => n10238, A2 => n10239, A3 => n10240, A4 => 
                           n10241, ZN => n7104);
   U6950 : AOI221_X1 port map( B1 => n19093, B2 => n10235, C1 => n19087, C2 => 
                           n10236, A => n10255, ZN => n10238);
   U6951 : AOI221_X1 port map( B1 => n19117, B2 => registers_15_20_port, C1 => 
                           n19111, C2 => registers_14_20_port, A => n10254, ZN 
                           => n10239);
   U6952 : NOR4_X1 port map( A1 => n10250, A2 => n10251, A3 => n10252, A4 => 
                           n10253, ZN => n10240);
   U6953 : NAND4_X1 port map( A1 => n10210, A2 => n10211, A3 => n10212, A4 => 
                           n10213, ZN => n7105);
   U6954 : AOI221_X1 port map( B1 => n19292, B2 => n10235, C1 => n19286, C2 => 
                           n10236, A => n10237, ZN => n10210);
   U6955 : NOR4_X1 port map( A1 => n10230, A2 => n10231, A3 => n10232, A4 => 
                           n10233, ZN => n10212);
   U6956 : AOI221_X1 port map( B1 => n19316, B2 => registers_15_20_port, C1 => 
                           n19310, C2 => registers_14_20_port, A => n10234, ZN 
                           => n10211);
   U6957 : NAND4_X1 port map( A1 => n10171, A2 => n10172, A3 => n10173, A4 => 
                           n10174, ZN => n7108);
   U6958 : AOI221_X1 port map( B1 => n19093, B2 => n10168, C1 => n19087, C2 => 
                           n10169, A => n10188, ZN => n10171);
   U6959 : AOI221_X1 port map( B1 => n19117, B2 => registers_15_21_port, C1 => 
                           n19111, C2 => registers_14_21_port, A => n10187, ZN 
                           => n10172);
   U6960 : NOR4_X1 port map( A1 => n10183, A2 => n10184, A3 => n10185, A4 => 
                           n10186, ZN => n10173);
   U6961 : NAND4_X1 port map( A1 => n10143, A2 => n10144, A3 => n10145, A4 => 
                           n10146, ZN => n7109);
   U6962 : AOI221_X1 port map( B1 => n19292, B2 => n10168, C1 => n19286, C2 => 
                           n10169, A => n10170, ZN => n10143);
   U6963 : NOR4_X1 port map( A1 => n10162, A2 => n10163, A3 => n10164, A4 => 
                           n10166, ZN => n10145);
   U6964 : AOI221_X1 port map( B1 => n19316, B2 => registers_15_21_port, C1 => 
                           n19310, C2 => registers_14_21_port, A => n10167, ZN 
                           => n10144);
   U6965 : NAND4_X1 port map( A1 => n10103, A2 => n10104, A3 => n10105, A4 => 
                           n10106, ZN => n7112);
   U6966 : AOI221_X1 port map( B1 => n19093, B2 => n10100, C1 => n19087, C2 => 
                           n10101, A => n10121, ZN => n10103);
   U6967 : AOI221_X1 port map( B1 => n19117, B2 => registers_15_22_port, C1 => 
                           n19111, C2 => registers_14_22_port, A => n10120, ZN 
                           => n10104);
   U6968 : NOR4_X1 port map( A1 => n10116, A2 => n10117, A3 => n10118, A4 => 
                           n10119, ZN => n10105);
   U6969 : NAND4_X1 port map( A1 => n10076, A2 => n10077, A3 => n10078, A4 => 
                           n10079, ZN => n7113);
   U6970 : AOI221_X1 port map( B1 => n19292, B2 => n10100, C1 => n19286, C2 => 
                           n10101, A => n10102, ZN => n10076);
   U6971 : NOR4_X1 port map( A1 => n10095, A2 => n10096, A3 => n10097, A4 => 
                           n10098, ZN => n10078);
   U6972 : AOI221_X1 port map( B1 => n19316, B2 => registers_15_22_port, C1 => 
                           n19310, C2 => registers_14_22_port, A => n10099, ZN 
                           => n10077);
   U6973 : NAND4_X1 port map( A1 => n10036, A2 => n10037, A3 => n10038, A4 => 
                           n10039, ZN => n7116);
   U6974 : AOI221_X1 port map( B1 => n19093, B2 => n10033, C1 => n19087, C2 => 
                           n10034, A => n10053, ZN => n10036);
   U6975 : AOI221_X1 port map( B1 => n19117, B2 => registers_15_23_port, C1 => 
                           n19111, C2 => registers_14_23_port, A => n10052, ZN 
                           => n10037);
   U6976 : NOR4_X1 port map( A1 => n10048, A2 => n10049, A3 => n10050, A4 => 
                           n10051, ZN => n10038);
   U6977 : NAND4_X1 port map( A1 => n10009, A2 => n10010, A3 => n10011, A4 => 
                           n10012, ZN => n7117);
   U6978 : AOI221_X1 port map( B1 => n19292, B2 => n10033, C1 => n19286, C2 => 
                           n10034, A => n10035, ZN => n10009);
   U6979 : NOR4_X1 port map( A1 => n10028, A2 => n10029, A3 => n10030, A4 => 
                           n10031, ZN => n10011);
   U6980 : AOI221_X1 port map( B1 => n19316, B2 => registers_15_23_port, C1 => 
                           n19310, C2 => registers_14_23_port, A => n10032, ZN 
                           => n10010);
   U6981 : NAND4_X1 port map( A1 => n9969, A2 => n9970, A3 => n9971, A4 => 
                           n9972, ZN => n7120);
   U6982 : AOI221_X1 port map( B1 => n19094, B2 => n9966, C1 => n19088, C2 => 
                           n9967, A => n9986, ZN => n9969);
   U6983 : AOI221_X1 port map( B1 => n19118, B2 => registers_15_24_port, C1 => 
                           n19112, C2 => registers_14_24_port, A => n9985, ZN 
                           => n9970);
   U6984 : NOR4_X1 port map( A1 => n9981, A2 => n9982, A3 => n9983, A4 => n9984
                           , ZN => n9971);
   U6985 : NAND4_X1 port map( A1 => n9941, A2 => n9942, A3 => n9943, A4 => 
                           n9944, ZN => n7121);
   U6986 : AOI221_X1 port map( B1 => n19293, B2 => n9966, C1 => n19287, C2 => 
                           n9967, A => n9968, ZN => n9941);
   U6987 : NOR4_X1 port map( A1 => n9961, A2 => n9962, A3 => n9963, A4 => n9964
                           , ZN => n9943);
   U6988 : AOI221_X1 port map( B1 => n19317, B2 => registers_15_24_port, C1 => 
                           n19311, C2 => registers_14_24_port, A => n9965, ZN 
                           => n9942);
   U6989 : NAND4_X1 port map( A1 => n9902, A2 => n9903, A3 => n9904, A4 => 
                           n9905, ZN => n7124);
   U6990 : AOI221_X1 port map( B1 => n19094, B2 => n9898, C1 => n19088, C2 => 
                           n9899, A => n9919, ZN => n9902);
   U6991 : AOI221_X1 port map( B1 => n19118, B2 => registers_15_25_port, C1 => 
                           n19112, C2 => registers_14_25_port, A => n9918, ZN 
                           => n9903);
   U6992 : NOR4_X1 port map( A1 => n9914, A2 => n9915, A3 => n9916, A4 => n9917
                           , ZN => n9904);
   U6993 : NAND4_X1 port map( A1 => n9874, A2 => n9875, A3 => n9876, A4 => 
                           n9877, ZN => n7125);
   U6994 : AOI221_X1 port map( B1 => n19293, B2 => n9898, C1 => n19287, C2 => 
                           n9899, A => n9900, ZN => n9874);
   U6995 : NOR4_X1 port map( A1 => n9893, A2 => n9894, A3 => n9895, A4 => n9896
                           , ZN => n9876);
   U6996 : AOI221_X1 port map( B1 => n19317, B2 => registers_15_25_port, C1 => 
                           n19311, C2 => registers_14_25_port, A => n9897, ZN 
                           => n9875);
   U6997 : NAND4_X1 port map( A1 => n9834, A2 => n9835, A3 => n9836, A4 => 
                           n9837, ZN => n7128);
   U6998 : AOI221_X1 port map( B1 => n19094, B2 => n9831, C1 => n19088, C2 => 
                           n9832, A => n9852, ZN => n9834);
   U6999 : AOI221_X1 port map( B1 => n19118, B2 => registers_15_26_port, C1 => 
                           n19112, C2 => registers_14_26_port, A => n9851, ZN 
                           => n9835);
   U7000 : NOR4_X1 port map( A1 => n9846, A2 => n9847, A3 => n9849, A4 => n9850
                           , ZN => n9836);
   U7001 : NAND4_X1 port map( A1 => n9807, A2 => n9808, A3 => n9809, A4 => 
                           n9810, ZN => n7129);
   U7002 : AOI221_X1 port map( B1 => n19293, B2 => n9831, C1 => n19287, C2 => 
                           n9832, A => n9833, ZN => n9807);
   U7003 : NOR4_X1 port map( A1 => n9826, A2 => n9827, A3 => n9828, A4 => n9829
                           , ZN => n9809);
   U7004 : AOI221_X1 port map( B1 => n19317, B2 => registers_15_26_port, C1 => 
                           n19311, C2 => registers_14_26_port, A => n9830, ZN 
                           => n9808);
   U7005 : NAND4_X1 port map( A1 => n9767, A2 => n9768, A3 => n9769, A4 => 
                           n9770, ZN => n7132);
   U7006 : AOI221_X1 port map( B1 => n19094, B2 => n9764, C1 => n19088, C2 => 
                           n9765, A => n9784, ZN => n9767);
   U7007 : AOI221_X1 port map( B1 => n19118, B2 => registers_15_27_port, C1 => 
                           n19112, C2 => registers_14_27_port, A => n9783, ZN 
                           => n9768);
   U7008 : NOR4_X1 port map( A1 => n9779, A2 => n9780, A3 => n9781, A4 => n9782
                           , ZN => n9769);
   U7009 : NAND4_X1 port map( A1 => n9739, A2 => n9740, A3 => n9741, A4 => 
                           n9743, ZN => n7133);
   U7010 : AOI221_X1 port map( B1 => n19293, B2 => n9764, C1 => n19287, C2 => 
                           n9765, A => n9766, ZN => n9739);
   U7011 : NOR4_X1 port map( A1 => n9759, A2 => n9760, A3 => n9761, A4 => n9762
                           , ZN => n9741);
   U7012 : AOI221_X1 port map( B1 => n19317, B2 => registers_15_27_port, C1 => 
                           n19311, C2 => registers_14_27_port, A => n9763, ZN 
                           => n9740);
   U7013 : NAND4_X1 port map( A1 => n9700, A2 => n9701, A3 => n9702, A4 => 
                           n9703, ZN => n7136);
   U7014 : AOI221_X1 port map( B1 => n19094, B2 => n9697, C1 => n19088, C2 => 
                           n9698, A => n9717, ZN => n9700);
   U7015 : AOI221_X1 port map( B1 => n19118, B2 => registers_15_28_port, C1 => 
                           n19112, C2 => registers_14_28_port, A => n9716, ZN 
                           => n9701);
   U7016 : NOR4_X1 port map( A1 => n9712, A2 => n9713, A3 => n9714, A4 => n9715
                           , ZN => n9702);
   U7017 : NAND4_X1 port map( A1 => n9672, A2 => n9673, A3 => n9674, A4 => 
                           n9675, ZN => n7137);
   U7018 : AOI221_X1 port map( B1 => n19293, B2 => n9697, C1 => n19287, C2 => 
                           n9698, A => n9699, ZN => n9672);
   U7019 : NOR4_X1 port map( A1 => n9692, A2 => n9693, A3 => n9694, A4 => n9695
                           , ZN => n9674);
   U7020 : AOI221_X1 port map( B1 => n19317, B2 => registers_15_28_port, C1 => 
                           n19311, C2 => registers_14_28_port, A => n9696, ZN 
                           => n9673);
   U7021 : NAND4_X1 port map( A1 => n9632, A2 => n9633, A3 => n9634, A4 => 
                           n9635, ZN => n7140);
   U7022 : AOI221_X1 port map( B1 => n19094, B2 => n9629, C1 => n19088, C2 => 
                           n9630, A => n9650, ZN => n9632);
   U7023 : AOI221_X1 port map( B1 => n19118, B2 => registers_15_29_port, C1 => 
                           n19112, C2 => registers_14_29_port, A => n9649, ZN 
                           => n9633);
   U7024 : NOR4_X1 port map( A1 => n9645, A2 => n9646, A3 => n9647, A4 => n9648
                           , ZN => n9634);
   U7025 : NAND4_X1 port map( A1 => n9605, A2 => n9606, A3 => n9607, A4 => 
                           n9608, ZN => n7141);
   U7026 : AOI221_X1 port map( B1 => n19293, B2 => n9629, C1 => n19287, C2 => 
                           n9630, A => n9631, ZN => n9605);
   U7027 : NOR4_X1 port map( A1 => n9624, A2 => n9625, A3 => n9626, A4 => n9627
                           , ZN => n9607);
   U7028 : AOI221_X1 port map( B1 => n19317, B2 => registers_15_29_port, C1 => 
                           n19311, C2 => registers_14_29_port, A => n9628, ZN 
                           => n9606);
   U7029 : NAND4_X1 port map( A1 => n9565, A2 => n9566, A3 => n9567, A4 => 
                           n9568, ZN => n7144);
   U7030 : AOI221_X1 port map( B1 => n19094, B2 => n9562, C1 => n19088, C2 => 
                           n9563, A => n9582, ZN => n9565);
   U7031 : AOI221_X1 port map( B1 => n19118, B2 => registers_15_30_port, C1 => 
                           n19112, C2 => registers_14_30_port, A => n9581, ZN 
                           => n9566);
   U7032 : NOR4_X1 port map( A1 => n9577, A2 => n9578, A3 => n9579, A4 => n9580
                           , ZN => n9567);
   U7033 : NAND4_X1 port map( A1 => n9538, A2 => n9539, A3 => n9540, A4 => 
                           n9541, ZN => n7145);
   U7034 : AOI221_X1 port map( B1 => n19293, B2 => n9562, C1 => n19287, C2 => 
                           n9563, A => n9564, ZN => n9538);
   U7035 : NOR4_X1 port map( A1 => n9557, A2 => n9558, A3 => n9559, A4 => n9560
                           , ZN => n9540);
   U7036 : AOI221_X1 port map( B1 => n19317, B2 => registers_15_30_port, C1 => 
                           n19311, C2 => registers_14_30_port, A => n9561, ZN 
                           => n9539);
   U7037 : NAND4_X1 port map( A1 => n9498, A2 => n9499, A3 => n9500, A4 => 
                           n9501, ZN => n7148);
   U7038 : AOI221_X1 port map( B1 => n19094, B2 => n9495, C1 => n19088, C2 => 
                           n9496, A => n9515, ZN => n9498);
   U7039 : AOI221_X1 port map( B1 => n19118, B2 => registers_15_31_port, C1 => 
                           n19112, C2 => registers_14_31_port, A => n9514, ZN 
                           => n9499);
   U7040 : NOR4_X1 port map( A1 => n9510, A2 => n9511, A3 => n9512, A4 => n9513
                           , ZN => n9500);
   U7041 : NAND4_X1 port map( A1 => n9470, A2 => n9471, A3 => n9472, A4 => 
                           n9473, ZN => n7149);
   U7042 : AOI221_X1 port map( B1 => n19293, B2 => n9495, C1 => n19287, C2 => 
                           n9496, A => n9497, ZN => n9470);
   U7043 : NOR4_X1 port map( A1 => n9490, A2 => n9491, A3 => n9492, A4 => n9493
                           , ZN => n9472);
   U7044 : AOI221_X1 port map( B1 => n19317, B2 => registers_15_31_port, C1 => 
                           n19311, C2 => registers_14_31_port, A => n9494, ZN 
                           => n9471);
   U7045 : NAND4_X1 port map( A1 => n9431, A2 => n9432, A3 => n9433, A4 => 
                           n9434, ZN => n7152);
   U7046 : AOI221_X1 port map( B1 => n19094, B2 => n9428, C1 => n19088, C2 => 
                           n9429, A => n9448, ZN => n9431);
   U7047 : AOI221_X1 port map( B1 => n19118, B2 => registers_15_32_port, C1 => 
                           n19112, C2 => registers_14_32_port, A => n9447, ZN 
                           => n9432);
   U7048 : NOR4_X1 port map( A1 => n9443, A2 => n9444, A3 => n9445, A4 => n9446
                           , ZN => n9433);
   U7049 : NAND4_X1 port map( A1 => n9403, A2 => n9404, A3 => n9405, A4 => 
                           n9406, ZN => n7153);
   U7050 : AOI221_X1 port map( B1 => n19293, B2 => n9428, C1 => n19287, C2 => 
                           n9429, A => n9430, ZN => n9403);
   U7051 : NOR4_X1 port map( A1 => n9422, A2 => n9423, A3 => n9425, A4 => n9426
                           , ZN => n9405);
   U7052 : AOI221_X1 port map( B1 => n19317, B2 => registers_15_32_port, C1 => 
                           n19311, C2 => registers_14_32_port, A => n9427, ZN 
                           => n9404);
   U7053 : NAND4_X1 port map( A1 => n9363, A2 => n9364, A3 => n9365, A4 => 
                           n9366, ZN => n7156);
   U7054 : AOI221_X1 port map( B1 => n19094, B2 => n9360, C1 => n19088, C2 => 
                           n9361, A => n9381, ZN => n9363);
   U7055 : AOI221_X1 port map( B1 => n19118, B2 => registers_15_33_port, C1 => 
                           n19112, C2 => registers_14_33_port, A => n9380, ZN 
                           => n9364);
   U7056 : NOR4_X1 port map( A1 => n9376, A2 => n9377, A3 => n9378, A4 => n9379
                           , ZN => n9365);
   U7057 : NAND4_X1 port map( A1 => n9336, A2 => n9337, A3 => n9338, A4 => 
                           n9339, ZN => n7157);
   U7058 : AOI221_X1 port map( B1 => n19293, B2 => n9360, C1 => n19287, C2 => 
                           n9361, A => n9362, ZN => n9336);
   U7059 : NOR4_X1 port map( A1 => n9355, A2 => n9356, A3 => n9357, A4 => n9358
                           , ZN => n9338);
   U7060 : AOI221_X1 port map( B1 => n19317, B2 => registers_15_33_port, C1 => 
                           n19311, C2 => registers_14_33_port, A => n9359, ZN 
                           => n9337);
   U7061 : NAND4_X1 port map( A1 => n9296, A2 => n9297, A3 => n9298, A4 => 
                           n9299, ZN => n7160);
   U7062 : AOI221_X1 port map( B1 => n19094, B2 => n9293, C1 => n19088, C2 => 
                           n9294, A => n9313, ZN => n9296);
   U7063 : AOI221_X1 port map( B1 => n19118, B2 => registers_15_34_port, C1 => 
                           n19112, C2 => registers_14_34_port, A => n9312, ZN 
                           => n9297);
   U7064 : NOR4_X1 port map( A1 => n9308, A2 => n9309, A3 => n9310, A4 => n9311
                           , ZN => n9298);
   U7065 : NAND4_X1 port map( A1 => n9269, A2 => n9270, A3 => n9271, A4 => 
                           n9272, ZN => n7161);
   U7066 : AOI221_X1 port map( B1 => n19293, B2 => n9293, C1 => n19287, C2 => 
                           n9294, A => n9295, ZN => n9269);
   U7067 : NOR4_X1 port map( A1 => n9288, A2 => n9289, A3 => n9290, A4 => n9291
                           , ZN => n9271);
   U7068 : AOI221_X1 port map( B1 => n19317, B2 => registers_15_34_port, C1 => 
                           n19311, C2 => registers_14_34_port, A => n9292, ZN 
                           => n9270);
   U7069 : NAND4_X1 port map( A1 => n6989, A2 => n6990, A3 => n6991, A4 => 
                           n6992, ZN => n7164);
   U7070 : AOI221_X1 port map( B1 => n19094, B2 => n6986, C1 => n19088, C2 => 
                           n6987, A => n7006, ZN => n6989);
   U7071 : AOI221_X1 port map( B1 => n19118, B2 => registers_15_35_port, C1 => 
                           n19112, C2 => registers_14_35_port, A => n7005, ZN 
                           => n6990);
   U7072 : NOR4_X1 port map( A1 => n7001, A2 => n7002, A3 => n7003, A4 => n7004
                           , ZN => n6991);
   U7073 : NAND4_X1 port map( A1 => n6962, A2 => n6963, A3 => n6964, A4 => 
                           n6965, ZN => n7165);
   U7074 : AOI221_X1 port map( B1 => n19293, B2 => n6986, C1 => n19287, C2 => 
                           n6987, A => n6988, ZN => n6962);
   U7075 : NOR4_X1 port map( A1 => n6981, A2 => n6982, A3 => n6983, A4 => n6984
                           , ZN => n6964);
   U7076 : AOI221_X1 port map( B1 => n19317, B2 => registers_15_35_port, C1 => 
                           n19311, C2 => registers_14_35_port, A => n6985, ZN 
                           => n6963);
   U7077 : NAND4_X1 port map( A1 => n6922, A2 => n6923, A3 => n6924, A4 => 
                           n6925, ZN => n7168);
   U7078 : AOI221_X1 port map( B1 => n19095, B2 => n6919, C1 => n19089, C2 => 
                           n6920, A => n6939, ZN => n6922);
   U7079 : AOI221_X1 port map( B1 => n19119, B2 => registers_15_36_port, C1 => 
                           n19113, C2 => registers_14_36_port, A => n6938, ZN 
                           => n6923);
   U7080 : NOR4_X1 port map( A1 => n6934, A2 => n6935, A3 => n6936, A4 => n6937
                           , ZN => n6924);
   U7081 : NAND4_X1 port map( A1 => n6895, A2 => n6896, A3 => n6897, A4 => 
                           n6898, ZN => n7169);
   U7082 : AOI221_X1 port map( B1 => n19294, B2 => n6919, C1 => n19288, C2 => 
                           n6920, A => n6921, ZN => n6895);
   U7083 : NOR4_X1 port map( A1 => n6914, A2 => n6915, A3 => n6916, A4 => n6917
                           , ZN => n6897);
   U7084 : AOI221_X1 port map( B1 => n19318, B2 => registers_15_36_port, C1 => 
                           n19312, C2 => registers_14_36_port, A => n6918, ZN 
                           => n6896);
   U7085 : NAND4_X1 port map( A1 => n6855, A2 => n6856, A3 => n6857, A4 => 
                           n6858, ZN => n7172);
   U7086 : AOI221_X1 port map( B1 => n19095, B2 => n6852, C1 => n19089, C2 => 
                           n6853, A => n6873, ZN => n6855);
   U7087 : AOI221_X1 port map( B1 => n19119, B2 => registers_15_37_port, C1 => 
                           n19113, C2 => registers_14_37_port, A => n6872, ZN 
                           => n6856);
   U7088 : NOR4_X1 port map( A1 => n6868, A2 => n6869, A3 => n6870, A4 => n6871
                           , ZN => n6857);
   U7089 : NAND4_X1 port map( A1 => n6828, A2 => n6829, A3 => n6830, A4 => 
                           n6831, ZN => n7173);
   U7090 : AOI221_X1 port map( B1 => n19294, B2 => n6852, C1 => n19288, C2 => 
                           n6853, A => n6854, ZN => n6828);
   U7091 : NOR4_X1 port map( A1 => n6847, A2 => n6848, A3 => n6849, A4 => n6850
                           , ZN => n6830);
   U7092 : AOI221_X1 port map( B1 => n19318, B2 => registers_15_37_port, C1 => 
                           n19312, C2 => registers_14_37_port, A => n6851, ZN 
                           => n6829);
   U7093 : NAND4_X1 port map( A1 => n6788, A2 => n6789, A3 => n6790, A4 => 
                           n6791, ZN => n7176);
   U7094 : AOI221_X1 port map( B1 => n19095, B2 => n6785, C1 => n19089, C2 => 
                           n6786, A => n6806, ZN => n6788);
   U7095 : AOI221_X1 port map( B1 => n19119, B2 => registers_15_38_port, C1 => 
                           n19113, C2 => registers_14_38_port, A => n6805, ZN 
                           => n6789);
   U7096 : NOR4_X1 port map( A1 => n6800, A2 => n6801, A3 => n6803, A4 => n6804
                           , ZN => n6790);
   U7097 : NAND4_X1 port map( A1 => n6761, A2 => n6762, A3 => n6763, A4 => 
                           n6764, ZN => n7177);
   U7098 : AOI221_X1 port map( B1 => n19294, B2 => n6785, C1 => n19288, C2 => 
                           n6786, A => n6787, ZN => n6761);
   U7099 : NOR4_X1 port map( A1 => n6780, A2 => n6781, A3 => n6782, A4 => n6783
                           , ZN => n6763);
   U7100 : AOI221_X1 port map( B1 => n19318, B2 => registers_15_38_port, C1 => 
                           n19312, C2 => registers_14_38_port, A => n6784, ZN 
                           => n6762);
   U7101 : NAND4_X1 port map( A1 => n6721, A2 => n6722, A3 => n6723, A4 => 
                           n6724, ZN => n7180);
   U7102 : AOI221_X1 port map( B1 => n19095, B2 => n6718, C1 => n19089, C2 => 
                           n6719, A => n6738, ZN => n6721);
   U7103 : AOI221_X1 port map( B1 => n19119, B2 => registers_15_39_port, C1 => 
                           n19113, C2 => registers_14_39_port, A => n6737, ZN 
                           => n6722);
   U7104 : NOR4_X1 port map( A1 => n6733, A2 => n6734, A3 => n6735, A4 => n6736
                           , ZN => n6723);
   U7105 : NAND4_X1 port map( A1 => n6693, A2 => n6694, A3 => n6695, A4 => 
                           n6697, ZN => n7181);
   U7106 : AOI221_X1 port map( B1 => n19294, B2 => n6718, C1 => n19288, C2 => 
                           n6719, A => n6720, ZN => n6693);
   U7107 : NOR4_X1 port map( A1 => n6713, A2 => n6714, A3 => n6715, A4 => n6716
                           , ZN => n6695);
   U7108 : AOI221_X1 port map( B1 => n19318, B2 => registers_15_39_port, C1 => 
                           n19312, C2 => registers_14_39_port, A => n6717, ZN 
                           => n6694);
   U7109 : NAND4_X1 port map( A1 => n6654, A2 => n6655, A3 => n6656, A4 => 
                           n6657, ZN => n7184);
   U7110 : AOI221_X1 port map( B1 => n19095, B2 => n6651, C1 => n19089, C2 => 
                           n6652, A => n6671, ZN => n6654);
   U7111 : AOI221_X1 port map( B1 => n19119, B2 => registers_15_40_port, C1 => 
                           n19113, C2 => registers_14_40_port, A => n6670, ZN 
                           => n6655);
   U7112 : NOR4_X1 port map( A1 => n6666, A2 => n6667, A3 => n6668, A4 => n6669
                           , ZN => n6656);
   U7113 : NAND4_X1 port map( A1 => n6626, A2 => n6627, A3 => n6628, A4 => 
                           n6629, ZN => n7185);
   U7114 : AOI221_X1 port map( B1 => n19294, B2 => n6651, C1 => n19288, C2 => 
                           n6652, A => n6653, ZN => n6626);
   U7115 : NOR4_X1 port map( A1 => n6646, A2 => n6647, A3 => n6648, A4 => n6649
                           , ZN => n6628);
   U7116 : AOI221_X1 port map( B1 => n19318, B2 => registers_15_40_port, C1 => 
                           n19312, C2 => registers_14_40_port, A => n6650, ZN 
                           => n6627);
   U7117 : NAND4_X1 port map( A1 => n6587, A2 => n6588, A3 => n6589, A4 => 
                           n6590, ZN => n7188);
   U7118 : AOI221_X1 port map( B1 => n19095, B2 => n6584, C1 => n19089, C2 => 
                           n6585, A => n6604, ZN => n6587);
   U7119 : AOI221_X1 port map( B1 => n19119, B2 => registers_15_41_port, C1 => 
                           n19113, C2 => registers_14_41_port, A => n6603, ZN 
                           => n6588);
   U7120 : NOR4_X1 port map( A1 => n6599, A2 => n6600, A3 => n6601, A4 => n6602
                           , ZN => n6589);
   U7121 : NAND4_X1 port map( A1 => n6560, A2 => n6561, A3 => n6562, A4 => 
                           n6563, ZN => n7189);
   U7122 : AOI221_X1 port map( B1 => n19294, B2 => n6584, C1 => n19288, C2 => 
                           n6585, A => n6586, ZN => n6560);
   U7123 : NOR4_X1 port map( A1 => n6579, A2 => n6580, A3 => n6581, A4 => n6582
                           , ZN => n6562);
   U7124 : AOI221_X1 port map( B1 => n19318, B2 => registers_15_41_port, C1 => 
                           n19312, C2 => registers_14_41_port, A => n6583, ZN 
                           => n6561);
   U7125 : NAND4_X1 port map( A1 => n6521, A2 => n6522, A3 => n6523, A4 => 
                           n6524, ZN => n7192);
   U7126 : AOI221_X1 port map( B1 => n19095, B2 => n6518, C1 => n19089, C2 => 
                           n6519, A => n6538, ZN => n6521);
   U7127 : AOI221_X1 port map( B1 => n19119, B2 => registers_15_42_port, C1 => 
                           n19113, C2 => registers_14_42_port, A => n6537, ZN 
                           => n6522);
   U7128 : NOR4_X1 port map( A1 => n6533, A2 => n6534, A3 => n6535, A4 => n6536
                           , ZN => n6523);
   U7129 : NAND4_X1 port map( A1 => n6494, A2 => n6495, A3 => n6496, A4 => 
                           n6497, ZN => n7193);
   U7130 : AOI221_X1 port map( B1 => n19294, B2 => n6518, C1 => n19288, C2 => 
                           n6519, A => n6520, ZN => n6494);
   U7131 : NOR4_X1 port map( A1 => n6513, A2 => n6514, A3 => n6515, A4 => n6516
                           , ZN => n6496);
   U7132 : AOI221_X1 port map( B1 => n19318, B2 => registers_15_42_port, C1 => 
                           n19312, C2 => registers_14_42_port, A => n6517, ZN 
                           => n6495);
   U7133 : NAND4_X1 port map( A1 => n6455, A2 => n6456, A3 => n6457, A4 => 
                           n6458, ZN => n7196);
   U7134 : AOI221_X1 port map( B1 => n19095, B2 => n6452, C1 => n19089, C2 => 
                           n6453, A => n6472, ZN => n6455);
   U7135 : AOI221_X1 port map( B1 => n19119, B2 => registers_15_43_port, C1 => 
                           n19113, C2 => registers_14_43_port, A => n6471, ZN 
                           => n6456);
   U7136 : NOR4_X1 port map( A1 => n6467, A2 => n6468, A3 => n6469, A4 => n6470
                           , ZN => n6457);
   U7137 : NAND4_X1 port map( A1 => n6428, A2 => n6429, A3 => n6430, A4 => 
                           n6431, ZN => n7197);
   U7138 : AOI221_X1 port map( B1 => n19294, B2 => n6452, C1 => n19288, C2 => 
                           n6453, A => n6454, ZN => n6428);
   U7139 : NOR4_X1 port map( A1 => n6447, A2 => n6448, A3 => n6449, A4 => n6450
                           , ZN => n6430);
   U7140 : AOI221_X1 port map( B1 => n19318, B2 => registers_15_43_port, C1 => 
                           n19312, C2 => registers_14_43_port, A => n6451, ZN 
                           => n6429);
   U7141 : NAND4_X1 port map( A1 => n6389, A2 => n6390, A3 => n6391, A4 => 
                           n6392, ZN => n7200);
   U7142 : AOI221_X1 port map( B1 => n19095, B2 => n6386, C1 => n19089, C2 => 
                           n6387, A => n6406, ZN => n6389);
   U7143 : AOI221_X1 port map( B1 => n19119, B2 => registers_15_44_port, C1 => 
                           n19113, C2 => registers_14_44_port, A => n6405, ZN 
                           => n6390);
   U7144 : NOR4_X1 port map( A1 => n6401, A2 => n6402, A3 => n6403, A4 => n6404
                           , ZN => n6391);
   U7145 : NAND4_X1 port map( A1 => n6362, A2 => n6363, A3 => n6364, A4 => 
                           n6365, ZN => n7201);
   U7146 : AOI221_X1 port map( B1 => n19294, B2 => n6386, C1 => n19288, C2 => 
                           n6387, A => n6388, ZN => n6362);
   U7147 : NOR4_X1 port map( A1 => n6381, A2 => n6382, A3 => n6383, A4 => n6384
                           , ZN => n6364);
   U7148 : AOI221_X1 port map( B1 => n19318, B2 => registers_15_44_port, C1 => 
                           n19312, C2 => registers_14_44_port, A => n6385, ZN 
                           => n6363);
   U7149 : NAND4_X1 port map( A1 => n6323, A2 => n6324, A3 => n6325, A4 => 
                           n6326, ZN => n7204);
   U7150 : AOI221_X1 port map( B1 => n19095, B2 => n6320, C1 => n19089, C2 => 
                           n6321, A => n6340, ZN => n6323);
   U7151 : AOI221_X1 port map( B1 => n19119, B2 => registers_15_45_port, C1 => 
                           n19113, C2 => registers_14_45_port, A => n6339, ZN 
                           => n6324);
   U7152 : NOR4_X1 port map( A1 => n6335, A2 => n6336, A3 => n6337, A4 => n6338
                           , ZN => n6325);
   U7153 : NAND4_X1 port map( A1 => n6296, A2 => n6297, A3 => n6298, A4 => 
                           n6299, ZN => n7205);
   U7154 : AOI221_X1 port map( B1 => n19294, B2 => n6320, C1 => n19288, C2 => 
                           n6321, A => n6322, ZN => n6296);
   U7155 : NOR4_X1 port map( A1 => n6315, A2 => n6316, A3 => n6317, A4 => n6318
                           , ZN => n6298);
   U7156 : AOI221_X1 port map( B1 => n19318, B2 => registers_15_45_port, C1 => 
                           n19312, C2 => registers_14_45_port, A => n6319, ZN 
                           => n6297);
   U7157 : NAND4_X1 port map( A1 => n6257, A2 => n6258, A3 => n6259, A4 => 
                           n6260, ZN => n7208);
   U7158 : AOI221_X1 port map( B1 => n19095, B2 => n6254, C1 => n19089, C2 => 
                           n6255, A => n6274, ZN => n6257);
   U7159 : AOI221_X1 port map( B1 => n19119, B2 => registers_15_46_port, C1 => 
                           n19113, C2 => registers_14_46_port, A => n6273, ZN 
                           => n6258);
   U7160 : NOR4_X1 port map( A1 => n6269, A2 => n6270, A3 => n6271, A4 => n6272
                           , ZN => n6259);
   U7161 : NAND4_X1 port map( A1 => n6230, A2 => n6231, A3 => n6232, A4 => 
                           n6233, ZN => n7209);
   U7162 : AOI221_X1 port map( B1 => n19294, B2 => n6254, C1 => n19288, C2 => 
                           n6255, A => n6256, ZN => n6230);
   U7163 : NOR4_X1 port map( A1 => n6249, A2 => n6250, A3 => n6251, A4 => n6252
                           , ZN => n6232);
   U7164 : AOI221_X1 port map( B1 => n19318, B2 => registers_15_46_port, C1 => 
                           n19312, C2 => registers_14_46_port, A => n6253, ZN 
                           => n6231);
   U7165 : NAND4_X1 port map( A1 => n6191, A2 => n6192, A3 => n6193, A4 => 
                           n6194, ZN => n7212);
   U7166 : AOI221_X1 port map( B1 => n19095, B2 => n6188, C1 => n19089, C2 => 
                           n6189, A => n6208, ZN => n6191);
   U7167 : AOI221_X1 port map( B1 => n19119, B2 => registers_15_47_port, C1 => 
                           n19113, C2 => registers_14_47_port, A => n6207, ZN 
                           => n6192);
   U7168 : NOR4_X1 port map( A1 => n6203, A2 => n6204, A3 => n6205, A4 => n6206
                           , ZN => n6193);
   U7169 : NAND4_X1 port map( A1 => n6164, A2 => n6165, A3 => n6166, A4 => 
                           n6167, ZN => n7213);
   U7170 : AOI221_X1 port map( B1 => n19294, B2 => n6188, C1 => n19288, C2 => 
                           n6189, A => n6190, ZN => n6164);
   U7171 : NOR4_X1 port map( A1 => n6183, A2 => n6184, A3 => n6185, A4 => n6186
                           , ZN => n6166);
   U7172 : AOI221_X1 port map( B1 => n19318, B2 => registers_15_47_port, C1 => 
                           n19312, C2 => registers_14_47_port, A => n6187, ZN 
                           => n6165);
   U7173 : NAND4_X1 port map( A1 => n6125, A2 => n6126, A3 => n6127, A4 => 
                           n6128, ZN => n7216);
   U7174 : AOI221_X1 port map( B1 => n19096, B2 => n6122, C1 => n19090, C2 => 
                           n6123, A => n6142, ZN => n6125);
   U7175 : AOI221_X1 port map( B1 => n19120, B2 => registers_15_48_port, C1 => 
                           n19114, C2 => registers_14_48_port, A => n6141, ZN 
                           => n6126);
   U7176 : NOR4_X1 port map( A1 => n6137, A2 => n6138, A3 => n6139, A4 => n6140
                           , ZN => n6127);
   U7177 : NAND4_X1 port map( A1 => n6098, A2 => n6099, A3 => n6100, A4 => 
                           n6101, ZN => n7217);
   U7178 : AOI221_X1 port map( B1 => n19295, B2 => n6122, C1 => n19289, C2 => 
                           n6123, A => n6124, ZN => n6098);
   U7179 : NOR4_X1 port map( A1 => n6117, A2 => n6118, A3 => n6119, A4 => n6120
                           , ZN => n6100);
   U7180 : AOI221_X1 port map( B1 => n19319, B2 => registers_15_48_port, C1 => 
                           n19313, C2 => registers_14_48_port, A => n6121, ZN 
                           => n6099);
   U7181 : NAND4_X1 port map( A1 => n6059, A2 => n6060, A3 => n6061, A4 => 
                           n6062, ZN => n7220);
   U7182 : AOI221_X1 port map( B1 => n19096, B2 => n6056, C1 => n19090, C2 => 
                           n6057, A => n6076, ZN => n6059);
   U7183 : AOI221_X1 port map( B1 => n19120, B2 => registers_15_49_port, C1 => 
                           n19114, C2 => registers_14_49_port, A => n6075, ZN 
                           => n6060);
   U7184 : NOR4_X1 port map( A1 => n6071, A2 => n6072, A3 => n6073, A4 => n6074
                           , ZN => n6061);
   U7185 : NAND4_X1 port map( A1 => n6030, A2 => n6031, A3 => n6032, A4 => 
                           n6034, ZN => n7221);
   U7186 : AOI221_X1 port map( B1 => n19295, B2 => n6056, C1 => n19289, C2 => 
                           n6057, A => n6058, ZN => n6030);
   U7187 : NOR4_X1 port map( A1 => n6051, A2 => n6052, A3 => n6053, A4 => n6054
                           , ZN => n6032);
   U7188 : AOI221_X1 port map( B1 => n19319, B2 => registers_15_49_port, C1 => 
                           n19313, C2 => registers_14_49_port, A => n6055, ZN 
                           => n6031);
   U7189 : NAND4_X1 port map( A1 => n5991, A2 => n5992, A3 => n5993, A4 => 
                           n5994, ZN => n7224);
   U7190 : AOI221_X1 port map( B1 => n19096, B2 => n5988, C1 => n19090, C2 => 
                           n5989, A => n6008, ZN => n5991);
   U7191 : AOI221_X1 port map( B1 => n19120, B2 => registers_15_50_port, C1 => 
                           n19114, C2 => registers_14_50_port, A => n6007, ZN 
                           => n5992);
   U7192 : NOR4_X1 port map( A1 => n6003, A2 => n6004, A3 => n6005, A4 => n6006
                           , ZN => n5993);
   U7193 : NAND4_X1 port map( A1 => n5962, A2 => n5963, A3 => n5964, A4 => 
                           n5965, ZN => n7225);
   U7194 : AOI221_X1 port map( B1 => n19295, B2 => n5988, C1 => n19289, C2 => 
                           n5989, A => n5990, ZN => n5962);
   U7195 : NOR4_X1 port map( A1 => n5983, A2 => n5984, A3 => n5985, A4 => n5986
                           , ZN => n5964);
   U7196 : AOI221_X1 port map( B1 => n19319, B2 => registers_15_50_port, C1 => 
                           n19313, C2 => registers_14_50_port, A => n5987, ZN 
                           => n5963);
   U7197 : NAND4_X1 port map( A1 => n5923, A2 => n5924, A3 => n5925, A4 => 
                           n5926, ZN => n7228);
   U7198 : AOI221_X1 port map( B1 => n19096, B2 => n5920, C1 => n19090, C2 => 
                           n5921, A => n5940, ZN => n5923);
   U7199 : AOI221_X1 port map( B1 => n19120, B2 => registers_15_51_port, C1 => 
                           n19114, C2 => registers_14_51_port, A => n5939, ZN 
                           => n5924);
   U7200 : NOR4_X1 port map( A1 => n5935, A2 => n5936, A3 => n5937, A4 => n5938
                           , ZN => n5925);
   U7201 : NAND4_X1 port map( A1 => n5895, A2 => n5896, A3 => n5897, A4 => 
                           n5898, ZN => n7229);
   U7202 : AOI221_X1 port map( B1 => n19295, B2 => n5920, C1 => n19289, C2 => 
                           n5921, A => n5922, ZN => n5895);
   U7203 : NOR4_X1 port map( A1 => n5915, A2 => n5916, A3 => n5917, A4 => n5918
                           , ZN => n5897);
   U7204 : AOI221_X1 port map( B1 => n19319, B2 => registers_15_51_port, C1 => 
                           n19313, C2 => registers_14_51_port, A => n5919, ZN 
                           => n5896);
   U7205 : NAND4_X1 port map( A1 => n5856, A2 => n5857, A3 => n5858, A4 => 
                           n5859, ZN => n7232);
   U7206 : AOI221_X1 port map( B1 => n19096, B2 => n5853, C1 => n19090, C2 => 
                           n5854, A => n5873, ZN => n5856);
   U7207 : AOI221_X1 port map( B1 => n19120, B2 => registers_15_52_port, C1 => 
                           n19114, C2 => registers_14_52_port, A => n5872, ZN 
                           => n5857);
   U7208 : NOR4_X1 port map( A1 => n5868, A2 => n5869, A3 => n5870, A4 => n5871
                           , ZN => n5858);
   U7209 : NAND4_X1 port map( A1 => n5828, A2 => n5829, A3 => n5830, A4 => 
                           n5831, ZN => n7233);
   U7210 : AOI221_X1 port map( B1 => n19295, B2 => n5853, C1 => n19289, C2 => 
                           n5854, A => n5855, ZN => n5828);
   U7211 : NOR4_X1 port map( A1 => n5848, A2 => n5849, A3 => n5850, A4 => n5851
                           , ZN => n5830);
   U7212 : AOI221_X1 port map( B1 => n19319, B2 => registers_15_52_port, C1 => 
                           n19313, C2 => registers_14_52_port, A => n5852, ZN 
                           => n5829);
   U7213 : NAND4_X1 port map( A1 => n5789, A2 => n5790, A3 => n5791, A4 => 
                           n5792, ZN => n7236);
   U7214 : AOI221_X1 port map( B1 => n19096, B2 => n5786, C1 => n19090, C2 => 
                           n5787, A => n5806, ZN => n5789);
   U7215 : AOI221_X1 port map( B1 => n19120, B2 => registers_15_53_port, C1 => 
                           n19114, C2 => registers_14_53_port, A => n5805, ZN 
                           => n5790);
   U7216 : NOR4_X1 port map( A1 => n5801, A2 => n5802, A3 => n5803, A4 => n5804
                           , ZN => n5791);
   U7217 : NAND4_X1 port map( A1 => n5756, A2 => n5757, A3 => n5758, A4 => 
                           n5759, ZN => n7237);
   U7218 : AOI221_X1 port map( B1 => n19295, B2 => n5786, C1 => n19289, C2 => 
                           n5787, A => n5788, ZN => n5756);
   U7219 : NOR4_X1 port map( A1 => n5781, A2 => n5782, A3 => n5783, A4 => n5784
                           , ZN => n5758);
   U7220 : AOI221_X1 port map( B1 => n19319, B2 => registers_15_53_port, C1 => 
                           n19313, C2 => registers_14_53_port, A => n5785, ZN 
                           => n5757);
   U7221 : NAND4_X1 port map( A1 => n5717, A2 => n5718, A3 => n5719, A4 => 
                           n5720, ZN => n7240);
   U7222 : AOI221_X1 port map( B1 => n19096, B2 => n5714, C1 => n19090, C2 => 
                           n5715, A => n5734, ZN => n5717);
   U7223 : AOI221_X1 port map( B1 => n19120, B2 => registers_15_54_port, C1 => 
                           n19114, C2 => registers_14_54_port, A => n5733, ZN 
                           => n5718);
   U7224 : NOR4_X1 port map( A1 => n5729, A2 => n5730, A3 => n5731, A4 => n5732
                           , ZN => n5719);
   U7225 : NAND4_X1 port map( A1 => n5686, A2 => n5687, A3 => n5688, A4 => 
                           n5689, ZN => n7241);
   U7226 : AOI221_X1 port map( B1 => n19295, B2 => n5714, C1 => n19289, C2 => 
                           n5715, A => n5716, ZN => n5686);
   U7227 : NOR4_X1 port map( A1 => n5709, A2 => n5710, A3 => n5711, A4 => n5712
                           , ZN => n5688);
   U7228 : AOI221_X1 port map( B1 => n19319, B2 => registers_15_54_port, C1 => 
                           n19313, C2 => registers_14_54_port, A => n5713, ZN 
                           => n5687);
   U7229 : NAND4_X1 port map( A1 => n5647, A2 => n5648, A3 => n5649, A4 => 
                           n5650, ZN => n7244);
   U7230 : AOI221_X1 port map( B1 => n19096, B2 => n5644, C1 => n19090, C2 => 
                           n5645, A => n5664, ZN => n5647);
   U7231 : AOI221_X1 port map( B1 => n19120, B2 => registers_15_55_port, C1 => 
                           n19114, C2 => registers_14_55_port, A => n5663, ZN 
                           => n5648);
   U7232 : NOR4_X1 port map( A1 => n5659, A2 => n5660, A3 => n5661, A4 => n5662
                           , ZN => n5649);
   U7233 : NAND4_X1 port map( A1 => n5618, A2 => n5619, A3 => n5620, A4 => 
                           n5621, ZN => n7245);
   U7234 : AOI221_X1 port map( B1 => n19295, B2 => n5644, C1 => n19289, C2 => 
                           n5645, A => n5646, ZN => n5618);
   U7235 : NOR4_X1 port map( A1 => n5639, A2 => n5640, A3 => n5641, A4 => n5642
                           , ZN => n5620);
   U7236 : AOI221_X1 port map( B1 => n19319, B2 => registers_15_55_port, C1 => 
                           n19313, C2 => registers_14_55_port, A => n5643, ZN 
                           => n5619);
   U7237 : NAND4_X1 port map( A1 => n5579, A2 => n5580, A3 => n5581, A4 => 
                           n5582, ZN => n7248);
   U7238 : AOI221_X1 port map( B1 => n19096, B2 => n5576, C1 => n19090, C2 => 
                           n5577, A => n5596, ZN => n5579);
   U7239 : AOI221_X1 port map( B1 => n19120, B2 => registers_15_56_port, C1 => 
                           n19114, C2 => registers_14_56_port, A => n5595, ZN 
                           => n5580);
   U7240 : NOR4_X1 port map( A1 => n5591, A2 => n5592, A3 => n5593, A4 => n5594
                           , ZN => n5581);
   U7241 : NAND4_X1 port map( A1 => n5549, A2 => n5550, A3 => n5551, A4 => 
                           n5552, ZN => n7249);
   U7242 : AOI221_X1 port map( B1 => n19295, B2 => n5576, C1 => n19289, C2 => 
                           n5577, A => n5578, ZN => n5549);
   U7243 : NOR4_X1 port map( A1 => n5571, A2 => n5572, A3 => n5573, A4 => n5574
                           , ZN => n5551);
   U7244 : AOI221_X1 port map( B1 => n19319, B2 => registers_15_56_port, C1 => 
                           n19313, C2 => registers_14_56_port, A => n5575, ZN 
                           => n5550);
   U7245 : NAND4_X1 port map( A1 => n5510, A2 => n5511, A3 => n5512, A4 => 
                           n5513, ZN => n7252);
   U7246 : AOI221_X1 port map( B1 => n19096, B2 => n5507, C1 => n19090, C2 => 
                           n5508, A => n5527, ZN => n5510);
   U7247 : AOI221_X1 port map( B1 => n19120, B2 => registers_15_57_port, C1 => 
                           n19114, C2 => registers_14_57_port, A => n5526, ZN 
                           => n5511);
   U7248 : NOR4_X1 port map( A1 => n5522, A2 => n5523, A3 => n5524, A4 => n5525
                           , ZN => n5512);
   U7249 : NAND4_X1 port map( A1 => n5480, A2 => n5481, A3 => n5482, A4 => 
                           n5483, ZN => n7253);
   U7250 : AOI221_X1 port map( B1 => n19295, B2 => n5507, C1 => n19289, C2 => 
                           n5508, A => n5509, ZN => n5480);
   U7251 : NOR4_X1 port map( A1 => n5502, A2 => n5503, A3 => n5504, A4 => n5505
                           , ZN => n5482);
   U7252 : AOI221_X1 port map( B1 => n19319, B2 => registers_15_57_port, C1 => 
                           n19313, C2 => registers_14_57_port, A => n5506, ZN 
                           => n5481);
   U7253 : NAND4_X1 port map( A1 => n5441, A2 => n5442, A3 => n5443, A4 => 
                           n5444, ZN => n7256);
   U7254 : AOI221_X1 port map( B1 => n19096, B2 => n5438, C1 => n19090, C2 => 
                           n5439, A => n5458, ZN => n5441);
   U7255 : AOI221_X1 port map( B1 => n19120, B2 => registers_15_58_port, C1 => 
                           n19114, C2 => registers_14_58_port, A => n5457, ZN 
                           => n5442);
   U7256 : NOR4_X1 port map( A1 => n5453, A2 => n5454, A3 => n5455, A4 => n5456
                           , ZN => n5443);
   U7257 : NAND4_X1 port map( A1 => n5412, A2 => n5413, A3 => n5414, A4 => 
                           n5415, ZN => n7257);
   U7258 : AOI221_X1 port map( B1 => n19295, B2 => n5438, C1 => n19289, C2 => 
                           n5439, A => n5440, ZN => n5412);
   U7259 : NOR4_X1 port map( A1 => n5433, A2 => n5434, A3 => n5435, A4 => n5436
                           , ZN => n5414);
   U7260 : AOI221_X1 port map( B1 => n19319, B2 => registers_15_58_port, C1 => 
                           n19313, C2 => registers_14_58_port, A => n5437, ZN 
                           => n5413);
   U7261 : NAND4_X1 port map( A1 => n5373, A2 => n5374, A3 => n5375, A4 => 
                           n5376, ZN => n7260);
   U7262 : AOI221_X1 port map( B1 => n19096, B2 => n5370, C1 => n19090, C2 => 
                           n5371, A => n5390, ZN => n5373);
   U7263 : AOI221_X1 port map( B1 => n19120, B2 => registers_15_59_port, C1 => 
                           n19114, C2 => registers_14_59_port, A => n5389, ZN 
                           => n5374);
   U7264 : NOR4_X1 port map( A1 => n5385, A2 => n5386, A3 => n5387, A4 => n5388
                           , ZN => n5375);
   U7265 : NAND4_X1 port map( A1 => n5342, A2 => n5343, A3 => n5344, A4 => 
                           n5345, ZN => n7261);
   U7266 : AOI221_X1 port map( B1 => n19295, B2 => n5370, C1 => n19289, C2 => 
                           n5371, A => n5372, ZN => n5342);
   U7267 : NOR4_X1 port map( A1 => n5365, A2 => n5366, A3 => n5367, A4 => n5368
                           , ZN => n5344);
   U7268 : AOI221_X1 port map( B1 => n19319, B2 => registers_15_59_port, C1 => 
                           n19313, C2 => registers_14_59_port, A => n5369, ZN 
                           => n5343);
   U7269 : NAND4_X1 port map( A1 => n5303, A2 => n5304, A3 => n5305, A4 => 
                           n5306, ZN => n7264);
   U7270 : AOI221_X1 port map( B1 => n19097, B2 => n5300, C1 => n19091, C2 => 
                           n5301, A => n5320, ZN => n5303);
   U7271 : AOI221_X1 port map( B1 => n19121, B2 => registers_15_60_port, C1 => 
                           n19115, C2 => registers_14_60_port, A => n5319, ZN 
                           => n5304);
   U7272 : NOR4_X1 port map( A1 => n5315, A2 => n5316, A3 => n5317, A4 => n5318
                           , ZN => n5305);
   U7273 : NAND4_X1 port map( A1 => n4857, A2 => n4922, A3 => n4923, A4 => 
                           n4988, ZN => n7265);
   U7274 : AOI221_X1 port map( B1 => n19296, B2 => n5300, C1 => n19290, C2 => 
                           n5301, A => n5302, ZN => n4857);
   U7275 : NOR4_X1 port map( A1 => n5295, A2 => n5296, A3 => n5297, A4 => n5298
                           , ZN => n4923);
   U7276 : AOI221_X1 port map( B1 => n19320, B2 => registers_15_60_port, C1 => 
                           n19314, C2 => registers_14_60_port, A => n5299, ZN 
                           => n4922);
   U7277 : NAND4_X1 port map( A1 => n4178, A2 => n4243, A3 => n4244, A4 => 
                           n4245, ZN => n7268);
   U7278 : AOI221_X1 port map( B1 => n19097, B2 => n4175, C1 => n19091, C2 => 
                           n4176, A => n4515, ZN => n4178);
   U7279 : AOI221_X1 port map( B1 => n19121, B2 => registers_15_61_port, C1 => 
                           n19115, C2 => registers_14_61_port, A => n4514, ZN 
                           => n4243);
   U7280 : NOR4_X1 port map( A1 => n4446, A2 => n4447, A3 => n4512, A4 => n4513
                           , ZN => n4244);
   U7281 : NAND4_X1 port map( A1 => n3639, A2 => n3640, A3 => n3705, A4 => 
                           n3706, ZN => n7269);
   U7282 : AOI221_X1 port map( B1 => n19296, B2 => n4175, C1 => n19290, C2 => 
                           n4176, A => n4177, ZN => n3639);
   U7283 : NOR4_X1 port map( A1 => n4106, A2 => n4107, A3 => n4108, A4 => n4109
                           , ZN => n3705);
   U7284 : AOI221_X1 port map( B1 => n19320, B2 => registers_15_61_port, C1 => 
                           n19314, C2 => registers_14_61_port, A => n4174, ZN 
                           => n3640);
   U7285 : NAND4_X1 port map( A1 => n3264, A2 => n3266, A3 => n3268, A4 => 
                           n3270, ZN => n7272);
   U7286 : AOI221_X1 port map( B1 => n19097, B2 => n3258, C1 => n19091, C2 => 
                           n3260, A => n3297, ZN => n3264);
   U7287 : AOI221_X1 port map( B1 => n19121, B2 => registers_15_62_port, C1 => 
                           n19115, C2 => registers_14_62_port, A => n3296, ZN 
                           => n3266);
   U7288 : NOR4_X1 port map( A1 => n3288, A2 => n3290, A3 => n3292, A4 => n3294
                           , ZN => n3268);
   U7289 : NAND4_X1 port map( A1 => n3210, A2 => n3212, A3 => n3214, A4 => 
                           n3216, ZN => n7273);
   U7290 : AOI221_X1 port map( B1 => n19296, B2 => n3258, C1 => n19290, C2 => 
                           n3260, A => n3262, ZN => n3210);
   U7291 : NOR4_X1 port map( A1 => n3248, A2 => n3250, A3 => n3252, A4 => n3254
                           , ZN => n3214);
   U7292 : AOI221_X1 port map( B1 => n19320, B2 => registers_15_62_port, C1 => 
                           n19314, C2 => registers_14_62_port, A => n3256, ZN 
                           => n3212);
   U7293 : NAND4_X1 port map( A1 => n3024, A2 => n3025, A3 => n3026, A4 => 
                           n3027, ZN => n7276);
   U7294 : AOI221_X1 port map( B1 => n19097, B2 => n3018, C1 => n19091, C2 => 
                           n3020, A => n3136, ZN => n3024);
   U7295 : AOI221_X1 port map( B1 => n19121, B2 => registers_15_63_port, C1 => 
                           n19115, C2 => registers_14_63_port, A => n3131, ZN 
                           => n3025);
   U7296 : NOR4_X1 port map( A1 => n3116, A2 => n3117, A3 => n3118, A4 => n3119
                           , ZN => n3026);
   U7297 : NAND4_X1 port map( A1 => n2772, A2 => n2773, A3 => n2774, A4 => 
                           n2775, ZN => n7277);
   U7298 : AOI221_X1 port map( B1 => n19296, B2 => n3018, C1 => n19290, C2 => 
                           n3020, A => n3021, ZN => n2772);
   U7299 : NOR4_X1 port map( A1 => n2999, A2 => n3000, A3 => n3001, A4 => n3002
                           , ZN => n2774);
   U7300 : AOI221_X1 port map( B1 => n19320, B2 => registers_15_63_port, C1 => 
                           n19314, C2 => registers_14_63_port, A => n3014, ZN 
                           => n2773);
   U7301 : NAND2_X1 port map( A1 => enable, A2 => n2092, ZN => n11557);
   U7302 : AND3_X1 port map( A1 => n11575, A2 => n20354, A3 => spill, ZN => 
                           n18902);
   U7303 : INV_X1 port map( A => count3(3), ZN => n11728);
   U7304 : NAND2_X1 port map( A1 => n11739, A2 => n11752, ZN => U3_U2_Z_3);
   U7305 : NAND2_X1 port map( A1 => n11739, A2 => n11751, ZN => U3_U6_Z_3);
   U7306 : NAND2_X1 port map( A1 => n11752, A2 => n11753, ZN => U3_U2_Z_1);
   U7307 : NAND2_X1 port map( A1 => n11751, A2 => n11753, ZN => U3_U6_Z_1);
   U7308 : NAND2_X1 port map( A1 => n11739, A2 => n11622, ZN => U3_U4_Z_3);
   U7309 : NAND2_X1 port map( A1 => n11622, A2 => n11753, ZN => U3_U4_Z_1);
   U7310 : OR3_X1 port map( A1 => n11671, A2 => count3(0), A3 => n11672, ZN => 
                           n11695);
   U7311 : AND3_X1 port map( A1 => n11671, A2 => n11672, A3 => count3(0), ZN =>
                           n11705);
   U7312 : INV_X1 port map( A => N92, ZN => n11749);
   U7313 : NOR2_X1 port map( A1 => U3_U2_Z_0, A2 => n11726, ZN => U3_U2_Z_4);
   U7314 : INV_X1 port map( A => N162, ZN => n11748);
   U7315 : NOR2_X1 port map( A1 => U3_U6_Z_0, A2 => n11726, ZN => U3_U6_Z_4);
   U7316 : INV_X1 port map( A => N127, ZN => n11623);
   U7317 : NOR2_X1 port map( A1 => U3_U4_Z_0, A2 => n11726, ZN => U3_U4_Z_4);
   U7318 : OR3_X1 port map( A1 => add_rd1(2), A2 => add_rd1(1), A3 => 
                           add_rd1(0), ZN => n11758);
   U7319 : OR3_X1 port map( A1 => add_wr(2), A2 => add_wr(1), A3 => add_wr(0), 
                           ZN => n11756);
   U7320 : INV_X1 port map( A => fill, ZN => n11575);
   U7321 : NOR2_X1 port map( A1 => n11575, A2 => reset, ZN => n2771);
   U7322 : NOR2_X1 port map( A1 => n2219, A2 => reset, ZN => n2770);
   U7323 : AOI22_X1 port map( A1 => datain(36), A2 => n19481, B1 => 
                           in_from_mem(36), B2 => n19475, ZN => n1660);
   U7324 : AOI22_X1 port map( A1 => datain(37), A2 => n19481, B1 => 
                           in_from_mem(37), B2 => n19475, ZN => n1659);
   U7325 : AOI22_X1 port map( A1 => datain(38), A2 => n19481, B1 => 
                           in_from_mem(38), B2 => n19475, ZN => n1658);
   U7326 : AOI22_X1 port map( A1 => datain(39), A2 => n19481, B1 => 
                           in_from_mem(39), B2 => n19475, ZN => n1657);
   U7327 : AOI22_X1 port map( A1 => datain(40), A2 => n19481, B1 => 
                           in_from_mem(40), B2 => n19475, ZN => n1656);
   U7328 : AOI22_X1 port map( A1 => datain(41), A2 => n19481, B1 => 
                           in_from_mem(41), B2 => n19475, ZN => n1655);
   U7329 : AOI22_X1 port map( A1 => datain(42), A2 => n19481, B1 => 
                           in_from_mem(42), B2 => n19475, ZN => n1654);
   U7330 : AOI22_X1 port map( A1 => datain(43), A2 => n19481, B1 => 
                           in_from_mem(43), B2 => n19475, ZN => n1653);
   U7331 : AOI22_X1 port map( A1 => datain(44), A2 => n19481, B1 => 
                           in_from_mem(44), B2 => n19475, ZN => n1652);
   U7332 : AOI22_X1 port map( A1 => datain(45), A2 => n19481, B1 => 
                           in_from_mem(45), B2 => n19475, ZN => n1651);
   U7333 : AOI22_X1 port map( A1 => datain(46), A2 => n19481, B1 => 
                           in_from_mem(46), B2 => n19475, ZN => n1650);
   U7334 : AOI22_X1 port map( A1 => datain(47), A2 => n19481, B1 => 
                           in_from_mem(47), B2 => n19475, ZN => n1649);
   U7335 : AOI22_X1 port map( A1 => datain(48), A2 => n19482, B1 => 
                           in_from_mem(48), B2 => n19476, ZN => n1648);
   U7336 : AOI22_X1 port map( A1 => datain(49), A2 => n19482, B1 => 
                           in_from_mem(49), B2 => n19476, ZN => n1647);
   U7337 : AOI22_X1 port map( A1 => datain(50), A2 => n19482, B1 => 
                           in_from_mem(50), B2 => n19476, ZN => n1646);
   U7338 : AOI22_X1 port map( A1 => datain(51), A2 => n19482, B1 => 
                           in_from_mem(51), B2 => n19476, ZN => n1645);
   U7339 : AOI22_X1 port map( A1 => datain(52), A2 => n19482, B1 => 
                           in_from_mem(52), B2 => n19476, ZN => n1644);
   U7340 : AOI22_X1 port map( A1 => datain(53), A2 => n19482, B1 => 
                           in_from_mem(53), B2 => n19476, ZN => n1643);
   U7341 : AOI22_X1 port map( A1 => datain(54), A2 => n19482, B1 => 
                           in_from_mem(54), B2 => n19476, ZN => n1642);
   U7342 : AOI22_X1 port map( A1 => datain(55), A2 => n19482, B1 => 
                           in_from_mem(55), B2 => n19476, ZN => n1641);
   U7343 : AOI22_X1 port map( A1 => datain(56), A2 => n19482, B1 => 
                           in_from_mem(56), B2 => n19476, ZN => n1640);
   U7344 : AOI22_X1 port map( A1 => datain(57), A2 => n19482, B1 => 
                           in_from_mem(57), B2 => n19476, ZN => n1639);
   U7345 : AOI22_X1 port map( A1 => datain(58), A2 => n19482, B1 => 
                           in_from_mem(58), B2 => n19476, ZN => n1638);
   U7346 : AOI22_X1 port map( A1 => datain(59), A2 => n19482, B1 => 
                           in_from_mem(59), B2 => n19476, ZN => n1637);
   U7347 : AOI22_X1 port map( A1 => datain(60), A2 => n19483, B1 => 
                           in_from_mem(60), B2 => n19477, ZN => n1636);
   U7348 : AOI22_X1 port map( A1 => datain(61), A2 => n19483, B1 => 
                           in_from_mem(61), B2 => n19477, ZN => n1635);
   U7349 : AOI22_X1 port map( A1 => datain(62), A2 => n19483, B1 => 
                           in_from_mem(62), B2 => n19477, ZN => n1634);
   U7350 : AOI22_X1 port map( A1 => datain(63), A2 => n19483, B1 => 
                           in_from_mem(63), B2 => n19477, ZN => n1631);
   U7351 : AOI22_X1 port map( A1 => datain(4), A2 => n19478, B1 => 
                           in_from_mem(4), B2 => n19472, ZN => n1692);
   U7352 : AOI22_X1 port map( A1 => datain(5), A2 => n19478, B1 => 
                           in_from_mem(5), B2 => n19472, ZN => n1691);
   U7353 : AOI22_X1 port map( A1 => datain(6), A2 => n19478, B1 => 
                           in_from_mem(6), B2 => n19472, ZN => n1690);
   U7354 : AOI22_X1 port map( A1 => datain(7), A2 => n19478, B1 => 
                           in_from_mem(7), B2 => n19472, ZN => n1689);
   U7355 : AOI22_X1 port map( A1 => datain(8), A2 => n19478, B1 => 
                           in_from_mem(8), B2 => n19472, ZN => n1688);
   U7356 : AOI22_X1 port map( A1 => datain(9), A2 => n19478, B1 => 
                           in_from_mem(9), B2 => n19472, ZN => n1687);
   U7357 : AOI22_X1 port map( A1 => datain(10), A2 => n19478, B1 => 
                           in_from_mem(10), B2 => n19472, ZN => n1686);
   U7358 : AOI22_X1 port map( A1 => datain(11), A2 => n19478, B1 => 
                           in_from_mem(11), B2 => n19472, ZN => n1685);
   U7359 : AOI22_X1 port map( A1 => datain(12), A2 => n19479, B1 => 
                           in_from_mem(12), B2 => n19473, ZN => n1684);
   U7360 : AOI22_X1 port map( A1 => datain(13), A2 => n19479, B1 => 
                           in_from_mem(13), B2 => n19473, ZN => n1683);
   U7361 : AOI22_X1 port map( A1 => datain(14), A2 => n19479, B1 => 
                           in_from_mem(14), B2 => n19473, ZN => n1682);
   U7362 : AOI22_X1 port map( A1 => datain(15), A2 => n19479, B1 => 
                           in_from_mem(15), B2 => n19473, ZN => n1681);
   U7363 : AOI22_X1 port map( A1 => datain(16), A2 => n19479, B1 => 
                           in_from_mem(16), B2 => n19473, ZN => n1680);
   U7364 : AOI22_X1 port map( A1 => datain(17), A2 => n19479, B1 => 
                           in_from_mem(17), B2 => n19473, ZN => n1679);
   U7365 : AOI22_X1 port map( A1 => datain(18), A2 => n19479, B1 => 
                           in_from_mem(18), B2 => n19473, ZN => n1678);
   U7366 : AOI22_X1 port map( A1 => datain(19), A2 => n19479, B1 => 
                           in_from_mem(19), B2 => n19473, ZN => n1677);
   U7367 : AOI22_X1 port map( A1 => datain(20), A2 => n19479, B1 => 
                           in_from_mem(20), B2 => n19473, ZN => n1676);
   U7368 : AOI22_X1 port map( A1 => datain(21), A2 => n19479, B1 => 
                           in_from_mem(21), B2 => n19473, ZN => n1675);
   U7369 : AOI22_X1 port map( A1 => datain(22), A2 => n19479, B1 => 
                           in_from_mem(22), B2 => n19473, ZN => n1674);
   U7370 : AOI22_X1 port map( A1 => datain(23), A2 => n19479, B1 => 
                           in_from_mem(23), B2 => n19473, ZN => n1673);
   U7371 : AOI22_X1 port map( A1 => datain(24), A2 => n19480, B1 => 
                           in_from_mem(24), B2 => n19474, ZN => n1672);
   U7372 : AOI22_X1 port map( A1 => datain(25), A2 => n19480, B1 => 
                           in_from_mem(25), B2 => n19474, ZN => n1671);
   U7373 : AOI22_X1 port map( A1 => datain(26), A2 => n19480, B1 => 
                           in_from_mem(26), B2 => n19474, ZN => n1670);
   U7375 : AOI22_X1 port map( A1 => datain(27), A2 => n19480, B1 => 
                           in_from_mem(27), B2 => n19474, ZN => n1669);
   U7376 : AOI22_X1 port map( A1 => datain(28), A2 => n19480, B1 => 
                           in_from_mem(28), B2 => n19474, ZN => n1668);
   U7377 : AOI22_X1 port map( A1 => datain(29), A2 => n19480, B1 => 
                           in_from_mem(29), B2 => n19474, ZN => n1667);
   U7378 : AOI22_X1 port map( A1 => datain(30), A2 => n19480, B1 => 
                           in_from_mem(30), B2 => n19474, ZN => n1666);
   U7379 : AOI22_X1 port map( A1 => datain(31), A2 => n19480, B1 => 
                           in_from_mem(31), B2 => n19474, ZN => n1665);
   U7380 : AOI22_X1 port map( A1 => datain(32), A2 => n19480, B1 => 
                           in_from_mem(32), B2 => n19474, ZN => n1664);
   U7381 : AOI22_X1 port map( A1 => datain(33), A2 => n19480, B1 => 
                           in_from_mem(33), B2 => n19474, ZN => n1663);
   U7382 : AOI22_X1 port map( A1 => datain(34), A2 => n19480, B1 => 
                           in_from_mem(34), B2 => n19474, ZN => n1662);
   U7383 : AOI22_X1 port map( A1 => datain(35), A2 => n19480, B1 => 
                           in_from_mem(35), B2 => n19474, ZN => n1661);
   U7384 : AOI22_X1 port map( A1 => datain(0), A2 => n19478, B1 => 
                           in_from_mem(0), B2 => n19472, ZN => n1696);
   U7385 : AOI22_X1 port map( A1 => datain(1), A2 => n19478, B1 => 
                           in_from_mem(1), B2 => n19472, ZN => n1695);
   U7386 : AOI22_X1 port map( A1 => datain(2), A2 => n19478, B1 => 
                           in_from_mem(2), B2 => n19472, ZN => n1694);
   U7387 : AOI22_X1 port map( A1 => datain(3), A2 => n19478, B1 => 
                           in_from_mem(3), B2 => n19472, ZN => n1693);
   U7388 : INV_X1 port map( A => count3(0), ZN => n1939);
   U7389 : NOR2_X1 port map( A1 => n11557, A2 => n11558, ZN => n2231);
   U7390 : INV_X1 port map( A => wr, ZN => n11558);
   U7391 : INV_X1 port map( A => reset, ZN => n1701);
   U7392 : INV_X1 port map( A => rd2, ZN => n11571);
   U7393 : NOR4_X1 port map( A1 => n6811, A2 => n6812, A3 => n6813, A4 => n6814
                           , ZN => n6810);
   U7394 : OAI221_X1 port map( B1 => n1825, B2 => n19053, C1 => n5282, C2 => 
                           n19047, A => n6815, ZN => n6813);
   U7395 : INV_X1 port map( A => n11747, ZN => n11562);
   U7396 : AOI221_X1 port map( B1 => n11654, B2 => n2764, C1 => N78, C2 => 
                           n2094, A => n11750, ZN => n11745);
   U7397 : AOI21_X1 port map( B1 => n11699, B2 => n11681, A => n2086, ZN => 
                           n11683);
   U7398 : OAI22_X1 port map( A1 => n4977, A2 => n18972, B1 => n5043, B2 => 
                           n18966, ZN => n10942);
   U7399 : OAI22_X1 port map( A1 => n4978, A2 => n18972, B1 => n5044, B2 => 
                           n18966, ZN => n11009);
   U7400 : OAI22_X1 port map( A1 => n4986, A2 => n18972, B1 => n5052, B2 => 
                           n18966, ZN => n11548);
   U7401 : OAI22_X1 port map( A1 => n4985, A2 => n18972, B1 => n5051, B2 => 
                           n18966, ZN => n11480);
   U7402 : OAI22_X1 port map( A1 => n4984, A2 => n18972, B1 => n5050, B2 => 
                           n18966, ZN => n11413);
   U7404 : OAI22_X1 port map( A1 => n4983, A2 => n18972, B1 => n5049, B2 => 
                           n18966, ZN => n11346);
   U7405 : OAI22_X1 port map( A1 => n4979, A2 => n18972, B1 => n5045, B2 => 
                           n18966, ZN => n11077);
   U7406 : OAI22_X1 port map( A1 => n4976, A2 => n18972, B1 => n5042, B2 => 
                           n18966, ZN => n10875);
   U7407 : OAI22_X1 port map( A1 => n4980, A2 => n18972, B1 => n5046, B2 => 
                           n18966, ZN => n11144);
   U7408 : OAI22_X1 port map( A1 => n4981, A2 => n18972, B1 => n5047, B2 => 
                           n18966, ZN => n11211);
   U7409 : OAI22_X1 port map( A1 => n4982, A2 => n18972, B1 => n5048, B2 => 
                           n18966, ZN => n11279);
   U7410 : OAI22_X1 port map( A1 => n4987, A2 => n18972, B1 => n5053, B2 => 
                           n18966, ZN => n11698);
   U7411 : OAI221_X1 port map( B1 => n1704, B2 => n2014, C1 => n1698, C2 => 
                           n2082, A => n20353, ZN => n2017);
   U7412 : OAI221_X1 port map( B1 => n1719, B2 => n2014, C1 => n1715, C2 => 
                           n2082, A => n20353, ZN => n2198);
   U7413 : OAI221_X1 port map( B1 => n1797, B2 => n2014, C1 => n1726, C2 => 
                           n2082, A => n20354, ZN => n2243);
   U7414 : OAI22_X1 port map( A1 => n11695, A2 => n11708, B1 => n2082, B2 => 
                           n11694, ZN => n11707);
   U7415 : OAI221_X1 port map( B1 => n1938, B2 => n2014, C1 => n1868, C2 => 
                           n2082, A => n20354, ZN => n2443);
   U7416 : NOR3_X1 port map( A1 => n11656, A2 => n11654, A3 => n11655, ZN => 
                           n11652);
   U7417 : AOI22_X1 port map( A1 => n11702, A2 => n2082, B1 => n11695, B2 => 
                           n11681, ZN => n11700);
   U7418 : NOR3_X1 port map( A1 => n11654, A2 => N78, A3 => n11656, ZN => 
                           n11645);
   U7419 : NOR3_X1 port map( A1 => n11563, A2 => n11656, A3 => n11655, ZN => 
                           n11642);
   U7420 : NOR3_X1 port map( A1 => n11656, A2 => N78, A3 => n11563, ZN => 
                           n11644);
   U7421 : INV_X1 port map( A => n11656, ZN => n11653);
   U7422 : NAND2_X1 port map( A1 => cwp(0), A2 => n11681, ZN => n11737);
   U7423 : NAND2_X1 port map( A1 => count3(1), A2 => cwp(0), ZN => n11731);
   U7424 : OAI22_X1 port map( A1 => n2092, A2 => n11728, B1 => n11656, B2 => 
                           n2219, ZN => n11747);
   U7425 : NAND2_X1 port map( A1 => cwp(1), A2 => cwp(0), ZN => n11726);
   U7426 : OAI221_X1 port map( B1 => n1709, B2 => n1938, C1 => n1712, C2 => 
                           n1868, A => n20353, ZN => n1945);
   U7427 : OAI221_X1 port map( B1 => n1699, B2 => n1938, C1 => n1705, C2 => 
                           n1868, A => n20353, ZN => n1873);
   U7428 : OAI221_X1 port map( B1 => n1697, B2 => n1868, C1 => n1699, C2 => 
                           n1869, A => n20352, ZN => n1867);
   U7429 : OAI221_X1 port map( B1 => n1708, B2 => n1868, C1 => n1709, C2 => 
                           n1869, A => n20353, ZN => n1942);
   U7430 : NAND2_X1 port map( A1 => n1940, A2 => n1947, ZN => n1709);
   U7431 : NAND2_X1 port map( A1 => n1940, A2 => N149, ZN => n1699);
   U7432 : OR3_X2 port map( A1 => n2091, A2 => n2092, A3 => n2093, ZN => n1698)
                           ;
   U7433 : NAND2_X1 port map( A1 => n11716, A2 => n2091, ZN => n2375);
   U7434 : NOR2_X1 port map( A1 => n2091, A2 => n11716, ZN => n2216);
   U7435 : XNOR2_X1 port map( A => n1940, B => n11574, ZN => n11566);
   U7436 : AOI21_X1 port map( B1 => n11731, B2 => n11732, A => n11733, ZN => 
                           n11729);
   U7437 : AOI21_X1 port map( B1 => n11734, B2 => n11735, A => count3(2), ZN =>
                           n11733);
   U7438 : OAI21_X1 port map( B1 => n11735, B2 => count3(2), A => n11734, ZN =>
                           n11740);
   U7459 : INV_X1 port map( A => n11744, ZN => n11559);
   U7464 : INV_X1 port map( A => n1940, ZN => n2764);
   U7469 : NAND2_X1 port map( A1 => n11732, A2 => n11622, ZN => U3_U4_Z_2);
   U7470 : NAND2_X1 port map( A1 => n11732, A2 => n11752, ZN => U3_U2_Z_2);
   U7471 : NAND2_X1 port map( A1 => n11732, A2 => n11751, ZN => U3_U6_Z_2);
   U7472 : INV_X1 port map( A => n11734, ZN => n11732);
   U7473 : OAI21_X1 port map( B1 => cwp(1), B2 => n11753, A => n11739, ZN => 
                           n11734);
   U7474 : OAI222_X1 port map( A1 => n11745, A2 => n2219, B1 => n11746, B2 => 
                           n2092, C1 => n2228, C2 => n11562, ZN => n11744);
   U7475 : BUF_X2 port map( A => n3170, Z => n18972);
   U7476 : CLKBUF_X1 port map( A => n3206, Z => n18908);
   U7477 : CLKBUF_X1 port map( A => n3202, Z => n18914);
   U7478 : CLKBUF_X1 port map( A => n3198, Z => n18923);
   U7479 : CLKBUF_X1 port map( A => n3196, Z => n18929);
   U7480 : CLKBUF_X1 port map( A => n3190, Z => n18935);
   U7481 : CLKBUF_X1 port map( A => n3186, Z => n18941);
   U7482 : CLKBUF_X1 port map( A => n3184, Z => n18947);
   U7483 : CLKBUF_X1 port map( A => n3180, Z => n18953);
   U7484 : CLKBUF_X1 port map( A => n3176, Z => n18959);
   U7485 : CLKBUF_X1 port map( A => n3174, Z => n18965);
   U7486 : CLKBUF_X1 port map( A => n3172, Z => n18971);
   U7487 : CLKBUF_X1 port map( A => n3170, Z => n18977);
   U7488 : CLKBUF_X1 port map( A => n3166, Z => n18983);
   U7489 : CLKBUF_X1 port map( A => n3165, Z => n18989);
   U7490 : CLKBUF_X1 port map( A => n3163, Z => n18995);
   U7491 : CLKBUF_X1 port map( A => n3161, Z => n19001);
   U7492 : CLKBUF_X1 port map( A => n3160, Z => n19007);
   U7493 : CLKBUF_X1 port map( A => n3159, Z => n19013);
   U7494 : CLKBUF_X1 port map( A => n3158, Z => n19019);
   U7495 : CLKBUF_X1 port map( A => n3156, Z => n19025);
   U7496 : CLKBUF_X1 port map( A => n3155, Z => n19031);
   U7497 : CLKBUF_X1 port map( A => n3154, Z => n19037);
   U7498 : CLKBUF_X1 port map( A => n3153, Z => n19043);
   U7499 : CLKBUF_X1 port map( A => n3151, Z => n19049);
   U7500 : CLKBUF_X1 port map( A => n3150, Z => n19055);
   U7501 : CLKBUF_X1 port map( A => n3149, Z => n19061);
   U7502 : CLKBUF_X1 port map( A => n3148, Z => n19067);
   U7503 : CLKBUF_X1 port map( A => n3147, Z => n19073);
   U7504 : CLKBUF_X1 port map( A => n3138, Z => n19079);
   U7505 : CLKBUF_X1 port map( A => n3137, Z => n19085);
   U7506 : CLKBUF_X1 port map( A => n3135, Z => n19091);
   U7507 : CLKBUF_X1 port map( A => n3134, Z => n19097);
   U7508 : CLKBUF_X1 port map( A => n3133, Z => n19103);
   U7509 : CLKBUF_X1 port map( A => n3132, Z => n19109);
   U7510 : CLKBUF_X1 port map( A => n3130, Z => n19115);
   U7511 : CLKBUF_X1 port map( A => n3129, Z => n19121);
   U7512 : CLKBUF_X1 port map( A => n3128, Z => n19127);
   U7513 : CLKBUF_X1 port map( A => n3127, Z => n19133);
   U7514 : CLKBUF_X1 port map( A => n3126, Z => n19139);
   U7515 : CLKBUF_X1 port map( A => n3125, Z => n19145);
   U7516 : CLKBUF_X1 port map( A => n3124, Z => n19151);
   U7517 : CLKBUF_X1 port map( A => n3123, Z => n19157);
   U7518 : CLKBUF_X1 port map( A => n3122, Z => n19163);
   U7519 : CLKBUF_X1 port map( A => n3120, Z => n19176);
   U7520 : CLKBUF_X1 port map( A => n3115, Z => n19182);
   U7521 : CLKBUF_X1 port map( A => n3114, Z => n19188);
   U7522 : CLKBUF_X1 port map( A => n3112, Z => n19194);
   U7523 : CLKBUF_X1 port map( A => n3111, Z => n19200);
   U7524 : CLKBUF_X1 port map( A => n3110, Z => n19206);
   U7525 : CLKBUF_X1 port map( A => n3109, Z => n19212);
   U7526 : CLKBUF_X1 port map( A => n3107, Z => n19218);
   U7527 : CLKBUF_X1 port map( A => n3106, Z => n19224);
   U7528 : CLKBUF_X1 port map( A => n3105, Z => n19230);
   U7529 : CLKBUF_X1 port map( A => n3104, Z => n19236);
   U7530 : CLKBUF_X1 port map( A => n3102, Z => n19242);
   U7531 : CLKBUF_X1 port map( A => n3037, Z => n19248);
   U7532 : CLKBUF_X1 port map( A => n3036, Z => n19254);
   U7533 : CLKBUF_X1 port map( A => n3035, Z => n19260);
   U7534 : CLKBUF_X1 port map( A => n3033, Z => n19266);
   U7535 : CLKBUF_X1 port map( A => n3032, Z => n19272);
   U7536 : CLKBUF_X1 port map( A => n3023, Z => n19278);
   U7537 : CLKBUF_X1 port map( A => n3022, Z => n19284);
   U7538 : CLKBUF_X1 port map( A => n3019, Z => n19290);
   U7539 : CLKBUF_X1 port map( A => n3017, Z => n19296);
   U7540 : CLKBUF_X1 port map( A => n3016, Z => n19302);
   U7541 : CLKBUF_X1 port map( A => n3015, Z => n19308);
   U7542 : CLKBUF_X1 port map( A => n3013, Z => n19314);
   U7543 : CLKBUF_X1 port map( A => n3012, Z => n19320);
   U7544 : CLKBUF_X1 port map( A => n3011, Z => n19326);
   U7545 : CLKBUF_X1 port map( A => n3010, Z => n19332);
   U7546 : CLKBUF_X1 port map( A => n3009, Z => n19338);
   U7547 : CLKBUF_X1 port map( A => n3008, Z => n19344);
   U7548 : CLKBUF_X1 port map( A => n3007, Z => n19350);
   U7549 : CLKBUF_X1 port map( A => n3006, Z => n19356);
   U7550 : CLKBUF_X1 port map( A => n3005, Z => n19362);
   U7551 : CLKBUF_X1 port map( A => n3003, Z => n19375);
   U7552 : CLKBUF_X1 port map( A => n2997, Z => n19381);
   U7553 : CLKBUF_X1 port map( A => n2995, Z => n19387);
   U7554 : CLKBUF_X1 port map( A => n2993, Z => n19393);
   U7555 : CLKBUF_X1 port map( A => n2992, Z => n19399);
   U7556 : CLKBUF_X1 port map( A => n2990, Z => n19405);
   U7557 : CLKBUF_X1 port map( A => n2988, Z => n19411);
   U7558 : CLKBUF_X1 port map( A => n2986, Z => n19417);
   U7559 : CLKBUF_X1 port map( A => n2985, Z => n19423);
   U7560 : CLKBUF_X1 port map( A => n2983, Z => n19429);
   U7561 : CLKBUF_X1 port map( A => n2982, Z => n19435);
   U7562 : CLKBUF_X1 port map( A => n2980, Z => n19441);
   U7563 : CLKBUF_X1 port map( A => n2979, Z => n19447);
   U7564 : CLKBUF_X1 port map( A => n2977, Z => n19453);
   U7565 : CLKBUF_X1 port map( A => n2783, Z => n19459);
   U7566 : CLKBUF_X1 port map( A => n2781, Z => n19465);
   U7567 : CLKBUF_X1 port map( A => n2780, Z => n19471);
   U7568 : CLKBUF_X1 port map( A => n2771, Z => n19477);
   U7569 : CLKBUF_X1 port map( A => n2770, Z => n19483);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_RF.all;

entity register_CU_A5_M8_N9_F4_B64_L32_T5_Y3 is

   port( clk, reset, call, ret : in std_logic;  spill, fill : out std_logic;  
         cwp : out std_logic_vector (1 downto 0);  count3 : out 
         std_logic_vector (3 downto 0));

end register_CU_A5_M8_N9_F4_B64_L32_T5_Y3;

architecture SYN_bhv of register_CU_A5_M8_N9_F4_B64_L32_T5_Y3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component register_CU_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_incdec_0
      port( A : in std_logic_vector (4 downto 0);  INC_DEC : in std_logic;  SUM
            : out std_logic_vector (4 downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal spill_port, fill_port, cwp_1_port, cwp_0_port, count3_3_port, 
      count3_2_port, count3_1_port, count3_0_port, swp_1_port, swp_0_port, 
      count_nested_4_port, count_nested_3_port, count_nested_2_port, 
      count_nested_1_port, count_nested_0_port, N192, N194, N196, N198, N200, 
      U3_U4_Z_0, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n111, n112, n114, n64, n65, n66, n67, n68, 
      n70, n71, n72, n73, n49, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n40, n41, n42, n44, n45, n46, n47, n48, n53, n54, n55, n56, 
      n57, n58, n59, n60, n61, n62, n63, n69, n74, n75, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93, n110, n113, n115
      , n116, n117, n119, n120, n121, n122 : std_logic;

begin
   spill <= spill_port;
   fill <= fill_port;
   cwp <= ( cwp_1_port, cwp_0_port );
   count3 <= ( count3_3_port, count3_2_port, count3_1_port, count3_0_port );
   
   temp_cwp_reg_0_inst : DFF_X1 port map( D => n108, CK => clk, Q => cwp_0_port
                           , QN => n70);
   count_nested_reg_3_inst : DFF_X1 port map( D => n107, CK => clk, Q => 
                           count_nested_3_port, QN => n68);
   must_fill_reg : DFF_X1 port map( D => n105, CK => clk, Q => fill_port, QN =>
                           n114);
   temp_count3_reg_2_inst : DFF_X1 port map( D => n104, CK => clk, Q => 
                           count3_2_port, QN => n111);
   temp_count3_reg_0_inst : DFF_X1 port map( D => n103, CK => clk, Q => 
                           count3_0_port, QN => n73);
   temp_count3_reg_1_inst : DFF_X1 port map( D => n102, CK => clk, Q => 
                           count3_1_port, QN => n72);
   temp_count3_reg_3_inst : DFF_X1 port map( D => n101, CK => clk, Q => 
                           count3_3_port, QN => n112);
   count_nested_reg_0_inst : DFF_X1 port map( D => n100, CK => clk, Q => 
                           count_nested_0_port, QN => n64);
   count_nested_reg_1_inst : DFF_X1 port map( D => n99, CK => clk, Q => 
                           count_nested_1_port, QN => n66);
   count_nested_reg_2_inst : DFF_X1 port map( D => n98, CK => clk, Q => 
                           count_nested_2_port, QN => n65);
   count_nested_reg_4_inst : DFF_X1 port map( D => n97, CK => clk, Q => 
                           count_nested_4_port, QN => n67);
   temp_cwp_reg_1_inst : DFF_X1 port map( D => n96, CK => clk, Q => cwp_1_port,
                           QN => n71);
   U76 : NAND3_X1 port map( A1 => n34, A2 => n35, A3 => n71, ZN => n33);
   U77 : NAND3_X1 port map( A1 => n44, A2 => n45, A3 => n114, ZN => n38);
   U78 : NAND3_X1 port map( A1 => cwp_0_port, A2 => cwp_1_port, A3 => n53, ZN 
                           => n48);
   U79 : NAND3_X1 port map( A1 => n37, A2 => n61, A3 => n63, ZN => n62);
   U80 : NAND3_X1 port map( A1 => n59, A2 => ret, A3 => n63, ZN => n78);
   U81 : XOR2_X1 port map( A => U3_U4_Z_0, B => cwp_0_port, Z => n35);
   U82 : NAND3_X1 port map( A1 => n111, A2 => count3_1_port, A3 => n90, ZN => 
                           n88);
   U83 : NAND3_X1 port map( A1 => n120, A2 => n122, A3 => call, ZN => U3_U4_Z_0
                           );
   r85 : register_CU_A5_M8_N9_F4_B64_L32_T5_Y3_DW01_incdec_0 port map( A(4) => 
                           count_nested_4_port, A(3) => count_nested_3_port, 
                           A(2) => count_nested_2_port, A(1) => 
                           count_nested_1_port, A(0) => count_nested_0_port, 
                           INC_DEC => U3_U4_Z_0, SUM(4) => N200, SUM(3) => N198
                           , SUM(2) => N196, SUM(1) => N194, SUM(0) => N192);
   flag_one_round_reg : DFF_X1 port map( D => n94, CK => clk, Q => n49, QN => 
                           n84);
   must_spill_reg : DFF_X1 port map( D => n109, CK => clk, Q => spill_port, QN 
                           => n56);
   swp_reg_0_inst : DFF_X1 port map( D => n106, CK => clk, Q => swp_0_port, QN 
                           => n61);
   swp_reg_1_inst : DFF_X1 port map( D => n95, CK => clk, Q => swp_1_port, QN 
                           => n40);
   U3 : INV_X1 port map( A => n92, ZN => n63);
   U4 : INV_X1 port map( A => n93, ZN => n119);
   U5 : INV_X1 port map( A => n28, ZN => n34);
   U6 : OAI211_X1 port map( C1 => n69, C2 => n74, A => n54, B => n45, ZN => n37
                           );
   U7 : NAND2_X1 port map( A1 => n69, A2 => n45, ZN => n27);
   U8 : INV_X1 port map( A => U3_U4_Z_0, ZN => n53);
   U9 : NAND2_X1 port map( A1 => n45, A2 => n27, ZN => n28);
   U10 : NOR2_X1 port map( A1 => n61, A2 => cwp_0_port, ZN => n83);
   U11 : OAI21_X1 port map( B1 => count3_1_port, B2 => n93, A => n113, ZN => 
                           n91);
   U12 : NAND2_X1 port map( A1 => n45, A2 => n86, ZN => n93);
   U13 : NAND2_X1 port map( A1 => n120, A2 => n45, ZN => n92);
   U14 : OAI21_X1 port map( B1 => n61, B2 => n37, A => n62, ZN => n106);
   U15 : INV_X1 port map( A => n90, ZN => n115);
   U16 : INV_X1 port map( A => n74, ZN => n59);
   U17 : INV_X1 port map( A => ret, ZN => n122);
   U18 : NOR2_X1 port map( A1 => fill_port, A2 => spill_port, ZN => n120);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n27, B1 => n28, B2 => n31, ZN => 
                           n97);
   U20 : INV_X1 port map( A => N200, ZN => n31);
   U21 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => n74);
   U22 : AOI221_X1 port map( B1 => n83, B2 => n53, C1 => n35, C2 => n61, A => 
                           n84, ZN => n79);
   U23 : AOI221_X1 port map( B1 => n42, B2 => n71, C1 => swp_1_port, C2 => n81,
                           A => n82, ZN => n80);
   U24 : NAND2_X1 port map( A1 => swp_0_port, A2 => U3_U4_Z_0, ZN => n46);
   U25 : NOR3_X1 port map( A1 => n63, A2 => n73, A3 => n93, ZN => n90);
   U26 : OAI22_X1 port map( A1 => n83, A2 => cwp_1_port, B1 => n71, B2 => n46, 
                           ZN => n81);
   U27 : AOI221_X1 port map( B1 => n37, B2 => n38, C1 => n40, C2 => n41, A => 
                           n42, ZN => n95);
   U28 : OAI21_X1 port map( B1 => swp_0_port, B2 => U3_U4_Z_0, A => n37, ZN => 
                           n41);
   U29 : AOI21_X1 port map( B1 => n73, B2 => n119, A => n63, ZN => n113);
   U30 : INV_X1 port map( A => reset, ZN => n45);
   U31 : AOI21_X1 port map( B1 => n120, B2 => ret, A => n53, ZN => n69);
   U32 : OAI211_X1 port map( C1 => swp_0_port, C2 => U3_U4_Z_0, A => n46, B => 
                           swp_1_port, ZN => n44);
   U33 : NOR3_X1 port map( A1 => n83, A2 => swp_1_port, A3 => n71, ZN => n82);
   U34 : NAND4_X1 port map( A1 => n73, A2 => n72, A3 => n111, A4 => 
                           count3_3_port, ZN => n86);
   U35 : OAI22_X1 port map( A1 => n65, A2 => n27, B1 => n28, B2 => n30, ZN => 
                           n98);
   U36 : INV_X1 port map( A => N196, ZN => n30);
   U37 : OAI22_X1 port map( A1 => n66, A2 => n27, B1 => n28, B2 => n29, ZN => 
                           n99);
   U38 : INV_X1 port map( A => N194, ZN => n29);
   U39 : OAI22_X1 port map( A1 => n64, A2 => n27, B1 => n28, B2 => n121, ZN => 
                           n100);
   U40 : INV_X1 port map( A => N192, ZN => n121);
   U41 : OAI22_X1 port map( A1 => n68, A2 => n27, B1 => n28, B2 => n60, ZN => 
                           n107);
   U42 : INV_X1 port map( A => N198, ZN => n60);
   U43 : OAI22_X1 port map( A1 => n70, A2 => n27, B1 => n28, B2 => cwp_0_port, 
                           ZN => n108);
   U44 : NOR2_X1 port map( A1 => n46, A2 => swp_1_port, ZN => n42);
   U45 : NOR2_X1 port map( A1 => n86, A2 => reset, ZN => n55);
   U46 : OAI22_X1 port map( A1 => n72, A2 => n113, B1 => count3_1_port, B2 => 
                           n115, ZN => n102);
   U47 : NAND4_X1 port map( A1 => n67, A2 => n66, A3 => n68, A4 => n75, ZN => 
                           n54);
   U48 : AND4_X1 port map( A1 => n56, A2 => fill_port, A3 => n64, A4 => n65, ZN
                           => n75);
   U49 : OAI21_X1 port map( B1 => n71, B2 => n32, A => n33, ZN => n96);
   U50 : INV_X1 port map( A => n36, ZN => n32);
   U51 : OAI21_X1 port map( B1 => n35, B2 => reset, A => n27, ZN => n36);
   U52 : AOI21_X1 port map( B1 => n47, B2 => n48, A => reset, ZN => n94);
   U53 : NAND2_X1 port map( A1 => n49, A2 => n54, ZN => n47);
   U54 : OAI21_X1 port map( B1 => n111, B2 => n87, A => n88, ZN => n104);
   U55 : INV_X1 port map( A => n91, ZN => n87);
   U56 : OAI21_X1 port map( B1 => n112, B2 => n116, A => n117, ZN => n101);
   U57 : AOI21_X1 port map( B1 => n119, B2 => n111, A => n91, ZN => n116);
   U58 : OR4_X1 port map( A1 => count3_3_port, A2 => n115, A3 => n111, A4 => 
                           n72, ZN => n117);
   U59 : OAI22_X1 port map( A1 => n73, A2 => n92, B1 => n93, B2 => n110, ZN => 
                           n103);
   U60 : NAND2_X1 port map( A1 => n73, A2 => n92, ZN => n110);
   U61 : OAI21_X1 port map( B1 => n55, B2 => n56, A => n57, ZN => n109);
   U62 : OAI211_X1 port map( C1 => n58, C2 => n59, A => n53, B => n45, ZN => 
                           n57);
   U63 : NOR3_X1 port map( A1 => n49, A2 => n71, A3 => n70, ZN => n58);
   U64 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => n105);
   U65 : OAI21_X1 port map( B1 => spill_port, B2 => n85, A => fill_port, ZN => 
                           n77);
   U66 : INV_X1 port map( A => n55, ZN => n85);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_RF.all;

entity windowed_RF is

   port( clk, reset, enable, call, ret, rd1, rd2, wr : in std_logic;  add_wr, 
         add_rd1, add_rd2 : in std_logic_vector (4 downto 0);  datain, 
         in_from_mem : in std_logic_vector (63 downto 0);  spill, fill : out 
         std_logic;  out_to_mem, out1, out2 : out std_logic_vector (63 downto 
         0));

end windowed_RF;

architecture SYN_struct of windowed_RF is

   component register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3
      port( clk, reset, enable, call, ret : in std_logic;  datain : in 
            std_logic_vector (63 downto 0);  rd1, rd2, wr : in std_logic;  
            add_wr, add_rd1, add_rd2 : in std_logic_vector (4 downto 0);  
            in_from_mem : in std_logic_vector (63 downto 0);  cwp : in 
            std_logic_vector (1 downto 0);  count3 : in std_logic_vector (3 
            downto 0);  spill, fill : in std_logic;  out_to_mem, out1, out2 : 
            out std_logic_vector (63 downto 0));
   end component;
   
   component register_CU_A5_M8_N9_F4_B64_L32_T5_Y3
      port( clk, reset, call, ret : in std_logic;  spill, fill : out std_logic;
            cwp : out std_logic_vector (1 downto 0);  count3 : out 
            std_logic_vector (3 downto 0));
   end component;
   
   signal spill_port, fill_port, temp_cwp_1_port, temp_cwp_0_port, 
      temp_count3_3_port, temp_count3_2_port, temp_count3_1_port, 
      temp_count3_0_port : std_logic;

begin
   spill <= spill_port;
   fill <= fill_port;
   
   Control_Unit : register_CU_A5_M8_N9_F4_B64_L32_T5_Y3 port map( clk => clk, 
                           reset => reset, call => call, ret => ret, spill => 
                           spill_port, fill => fill_port, cwp(1) => 
                           temp_cwp_1_port, cwp(0) => temp_cwp_0_port, 
                           count3(3) => temp_count3_3_port, count3(2) => 
                           temp_count3_2_port, count3(1) => temp_count3_1_port,
                           count3(0) => temp_count3_0_port);
   Register_File_and_addresses : register_file_w_A5_M8_N9_F4_B64_L32_T5_Y3 port
                           map( clk => clk, reset => reset, enable => enable, 
                           call => call, ret => ret, datain(63) => datain(63), 
                           datain(62) => datain(62), datain(61) => datain(61), 
                           datain(60) => datain(60), datain(59) => datain(59), 
                           datain(58) => datain(58), datain(57) => datain(57), 
                           datain(56) => datain(56), datain(55) => datain(55), 
                           datain(54) => datain(54), datain(53) => datain(53), 
                           datain(52) => datain(52), datain(51) => datain(51), 
                           datain(50) => datain(50), datain(49) => datain(49), 
                           datain(48) => datain(48), datain(47) => datain(47), 
                           datain(46) => datain(46), datain(45) => datain(45), 
                           datain(44) => datain(44), datain(43) => datain(43), 
                           datain(42) => datain(42), datain(41) => datain(41), 
                           datain(40) => datain(40), datain(39) => datain(39), 
                           datain(38) => datain(38), datain(37) => datain(37), 
                           datain(36) => datain(36), datain(35) => datain(35), 
                           datain(34) => datain(34), datain(33) => datain(33), 
                           datain(32) => datain(32), datain(31) => datain(31), 
                           datain(30) => datain(30), datain(29) => datain(29), 
                           datain(28) => datain(28), datain(27) => datain(27), 
                           datain(26) => datain(26), datain(25) => datain(25), 
                           datain(24) => datain(24), datain(23) => datain(23), 
                           datain(22) => datain(22), datain(21) => datain(21), 
                           datain(20) => datain(20), datain(19) => datain(19), 
                           datain(18) => datain(18), datain(17) => datain(17), 
                           datain(16) => datain(16), datain(15) => datain(15), 
                           datain(14) => datain(14), datain(13) => datain(13), 
                           datain(12) => datain(12), datain(11) => datain(11), 
                           datain(10) => datain(10), datain(9) => datain(9), 
                           datain(8) => datain(8), datain(7) => datain(7), 
                           datain(6) => datain(6), datain(5) => datain(5), 
                           datain(4) => datain(4), datain(3) => datain(3), 
                           datain(2) => datain(2), datain(1) => datain(1), 
                           datain(0) => datain(0), rd1 => rd1, rd2 => rd2, wr 
                           => wr, add_wr(4) => add_wr(4), add_wr(3) => 
                           add_wr(3), add_wr(2) => add_wr(2), add_wr(1) => 
                           add_wr(1), add_wr(0) => add_wr(0), add_rd1(4) => 
                           add_rd1(4), add_rd1(3) => add_rd1(3), add_rd1(2) => 
                           add_rd1(2), add_rd1(1) => add_rd1(1), add_rd1(0) => 
                           add_rd1(0), add_rd2(4) => add_rd2(4), add_rd2(3) => 
                           add_rd2(3), add_rd2(2) => add_rd2(2), add_rd2(1) => 
                           add_rd2(1), add_rd2(0) => add_rd2(0), 
                           in_from_mem(63) => in_from_mem(63), in_from_mem(62) 
                           => in_from_mem(62), in_from_mem(61) => 
                           in_from_mem(61), in_from_mem(60) => in_from_mem(60),
                           in_from_mem(59) => in_from_mem(59), in_from_mem(58) 
                           => in_from_mem(58), in_from_mem(57) => 
                           in_from_mem(57), in_from_mem(56) => in_from_mem(56),
                           in_from_mem(55) => in_from_mem(55), in_from_mem(54) 
                           => in_from_mem(54), in_from_mem(53) => 
                           in_from_mem(53), in_from_mem(52) => in_from_mem(52),
                           in_from_mem(51) => in_from_mem(51), in_from_mem(50) 
                           => in_from_mem(50), in_from_mem(49) => 
                           in_from_mem(49), in_from_mem(48) => in_from_mem(48),
                           in_from_mem(47) => in_from_mem(47), in_from_mem(46) 
                           => in_from_mem(46), in_from_mem(45) => 
                           in_from_mem(45), in_from_mem(44) => in_from_mem(44),
                           in_from_mem(43) => in_from_mem(43), in_from_mem(42) 
                           => in_from_mem(42), in_from_mem(41) => 
                           in_from_mem(41), in_from_mem(40) => in_from_mem(40),
                           in_from_mem(39) => in_from_mem(39), in_from_mem(38) 
                           => in_from_mem(38), in_from_mem(37) => 
                           in_from_mem(37), in_from_mem(36) => in_from_mem(36),
                           in_from_mem(35) => in_from_mem(35), in_from_mem(34) 
                           => in_from_mem(34), in_from_mem(33) => 
                           in_from_mem(33), in_from_mem(32) => in_from_mem(32),
                           in_from_mem(31) => in_from_mem(31), in_from_mem(30) 
                           => in_from_mem(30), in_from_mem(29) => 
                           in_from_mem(29), in_from_mem(28) => in_from_mem(28),
                           in_from_mem(27) => in_from_mem(27), in_from_mem(26) 
                           => in_from_mem(26), in_from_mem(25) => 
                           in_from_mem(25), in_from_mem(24) => in_from_mem(24),
                           in_from_mem(23) => in_from_mem(23), in_from_mem(22) 
                           => in_from_mem(22), in_from_mem(21) => 
                           in_from_mem(21), in_from_mem(20) => in_from_mem(20),
                           in_from_mem(19) => in_from_mem(19), in_from_mem(18) 
                           => in_from_mem(18), in_from_mem(17) => 
                           in_from_mem(17), in_from_mem(16) => in_from_mem(16),
                           in_from_mem(15) => in_from_mem(15), in_from_mem(14) 
                           => in_from_mem(14), in_from_mem(13) => 
                           in_from_mem(13), in_from_mem(12) => in_from_mem(12),
                           in_from_mem(11) => in_from_mem(11), in_from_mem(10) 
                           => in_from_mem(10), in_from_mem(9) => in_from_mem(9)
                           , in_from_mem(8) => in_from_mem(8), in_from_mem(7) 
                           => in_from_mem(7), in_from_mem(6) => in_from_mem(6),
                           in_from_mem(5) => in_from_mem(5), in_from_mem(4) => 
                           in_from_mem(4), in_from_mem(3) => in_from_mem(3), 
                           in_from_mem(2) => in_from_mem(2), in_from_mem(1) => 
                           in_from_mem(1), in_from_mem(0) => in_from_mem(0), 
                           cwp(1) => temp_cwp_1_port, cwp(0) => temp_cwp_0_port
                           , count3(3) => temp_count3_3_port, count3(2) => 
                           temp_count3_2_port, count3(1) => temp_count3_1_port,
                           count3(0) => temp_count3_0_port, spill => spill_port
                           , fill => fill_port, out_to_mem(63) => 
                           out_to_mem(63), out_to_mem(62) => out_to_mem(62), 
                           out_to_mem(61) => out_to_mem(61), out_to_mem(60) => 
                           out_to_mem(60), out_to_mem(59) => out_to_mem(59), 
                           out_to_mem(58) => out_to_mem(58), out_to_mem(57) => 
                           out_to_mem(57), out_to_mem(56) => out_to_mem(56), 
                           out_to_mem(55) => out_to_mem(55), out_to_mem(54) => 
                           out_to_mem(54), out_to_mem(53) => out_to_mem(53), 
                           out_to_mem(52) => out_to_mem(52), out_to_mem(51) => 
                           out_to_mem(51), out_to_mem(50) => out_to_mem(50), 
                           out_to_mem(49) => out_to_mem(49), out_to_mem(48) => 
                           out_to_mem(48), out_to_mem(47) => out_to_mem(47), 
                           out_to_mem(46) => out_to_mem(46), out_to_mem(45) => 
                           out_to_mem(45), out_to_mem(44) => out_to_mem(44), 
                           out_to_mem(43) => out_to_mem(43), out_to_mem(42) => 
                           out_to_mem(42), out_to_mem(41) => out_to_mem(41), 
                           out_to_mem(40) => out_to_mem(40), out_to_mem(39) => 
                           out_to_mem(39), out_to_mem(38) => out_to_mem(38), 
                           out_to_mem(37) => out_to_mem(37), out_to_mem(36) => 
                           out_to_mem(36), out_to_mem(35) => out_to_mem(35), 
                           out_to_mem(34) => out_to_mem(34), out_to_mem(33) => 
                           out_to_mem(33), out_to_mem(32) => out_to_mem(32), 
                           out_to_mem(31) => out_to_mem(31), out_to_mem(30) => 
                           out_to_mem(30), out_to_mem(29) => out_to_mem(29), 
                           out_to_mem(28) => out_to_mem(28), out_to_mem(27) => 
                           out_to_mem(27), out_to_mem(26) => out_to_mem(26), 
                           out_to_mem(25) => out_to_mem(25), out_to_mem(24) => 
                           out_to_mem(24), out_to_mem(23) => out_to_mem(23), 
                           out_to_mem(22) => out_to_mem(22), out_to_mem(21) => 
                           out_to_mem(21), out_to_mem(20) => out_to_mem(20), 
                           out_to_mem(19) => out_to_mem(19), out_to_mem(18) => 
                           out_to_mem(18), out_to_mem(17) => out_to_mem(17), 
                           out_to_mem(16) => out_to_mem(16), out_to_mem(15) => 
                           out_to_mem(15), out_to_mem(14) => out_to_mem(14), 
                           out_to_mem(13) => out_to_mem(13), out_to_mem(12) => 
                           out_to_mem(12), out_to_mem(11) => out_to_mem(11), 
                           out_to_mem(10) => out_to_mem(10), out_to_mem(9) => 
                           out_to_mem(9), out_to_mem(8) => out_to_mem(8), 
                           out_to_mem(7) => out_to_mem(7), out_to_mem(6) => 
                           out_to_mem(6), out_to_mem(5) => out_to_mem(5), 
                           out_to_mem(4) => out_to_mem(4), out_to_mem(3) => 
                           out_to_mem(3), out_to_mem(2) => out_to_mem(2), 
                           out_to_mem(1) => out_to_mem(1), out_to_mem(0) => 
                           out_to_mem(0), out1(63) => out1(63), out1(62) => 
                           out1(62), out1(61) => out1(61), out1(60) => out1(60)
                           , out1(59) => out1(59), out1(58) => out1(58), 
                           out1(57) => out1(57), out1(56) => out1(56), out1(55)
                           => out1(55), out1(54) => out1(54), out1(53) => 
                           out1(53), out1(52) => out1(52), out1(51) => out1(51)
                           , out1(50) => out1(50), out1(49) => out1(49), 
                           out1(48) => out1(48), out1(47) => out1(47), out1(46)
                           => out1(46), out1(45) => out1(45), out1(44) => 
                           out1(44), out1(43) => out1(43), out1(42) => out1(42)
                           , out1(41) => out1(41), out1(40) => out1(40), 
                           out1(39) => out1(39), out1(38) => out1(38), out1(37)
                           => out1(37), out1(36) => out1(36), out1(35) => 
                           out1(35), out1(34) => out1(34), out1(33) => out1(33)
                           , out1(32) => out1(32), out1(31) => out1(31), 
                           out1(30) => out1(30), out1(29) => out1(29), out1(28)
                           => out1(28), out1(27) => out1(27), out1(26) => 
                           out1(26), out1(25) => out1(25), out1(24) => out1(24)
                           , out1(23) => out1(23), out1(22) => out1(22), 
                           out1(21) => out1(21), out1(20) => out1(20), out1(19)
                           => out1(19), out1(18) => out1(18), out1(17) => 
                           out1(17), out1(16) => out1(16), out1(15) => out1(15)
                           , out1(14) => out1(14), out1(13) => out1(13), 
                           out1(12) => out1(12), out1(11) => out1(11), out1(10)
                           => out1(10), out1(9) => out1(9), out1(8) => out1(8),
                           out1(7) => out1(7), out1(6) => out1(6), out1(5) => 
                           out1(5), out1(4) => out1(4), out1(3) => out1(3), 
                           out1(2) => out1(2), out1(1) => out1(1), out1(0) => 
                           out1(0), out2(63) => out2(63), out2(62) => out2(62),
                           out2(61) => out2(61), out2(60) => out2(60), out2(59)
                           => out2(59), out2(58) => out2(58), out2(57) => 
                           out2(57), out2(56) => out2(56), out2(55) => out2(55)
                           , out2(54) => out2(54), out2(53) => out2(53), 
                           out2(52) => out2(52), out2(51) => out2(51), out2(50)
                           => out2(50), out2(49) => out2(49), out2(48) => 
                           out2(48), out2(47) => out2(47), out2(46) => out2(46)
                           , out2(45) => out2(45), out2(44) => out2(44), 
                           out2(43) => out2(43), out2(42) => out2(42), out2(41)
                           => out2(41), out2(40) => out2(40), out2(39) => 
                           out2(39), out2(38) => out2(38), out2(37) => out2(37)
                           , out2(36) => out2(36), out2(35) => out2(35), 
                           out2(34) => out2(34), out2(33) => out2(33), out2(32)
                           => out2(32), out2(31) => out2(31), out2(30) => 
                           out2(30), out2(29) => out2(29), out2(28) => out2(28)
                           , out2(27) => out2(27), out2(26) => out2(26), 
                           out2(25) => out2(25), out2(24) => out2(24), out2(23)
                           => out2(23), out2(22) => out2(22), out2(21) => 
                           out2(21), out2(20) => out2(20), out2(19) => out2(19)
                           , out2(18) => out2(18), out2(17) => out2(17), 
                           out2(16) => out2(16), out2(15) => out2(15), out2(14)
                           => out2(14), out2(13) => out2(13), out2(12) => 
                           out2(12), out2(11) => out2(11), out2(10) => out2(10)
                           , out2(9) => out2(9), out2(8) => out2(8), out2(7) =>
                           out2(7), out2(6) => out2(6), out2(5) => out2(5), 
                           out2(4) => out2(4), out2(3) => out2(3), out2(2) => 
                           out2(2), out2(1) => out2(1), out2(0) => out2(0));

end SYN_struct;
