package CONSTANTS is


	constant num_bit : integer := 32;
	constant global 	: integer := 4; 
	constant win 		: integer := 4;                     --- 32 X 36
	constant dimension_in_local_out : integer := 4;
	
	constant max_nested_calls : integer := 32;
	
	
end CONSTANTS;
