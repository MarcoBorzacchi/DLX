package CONSTANTS is

	constant NumBit : integer := 32;
	constant numBit_block : integer := 4;
	constant n_blocks : integer := 8;
 	
end CONSTANTS;
